module RS(
  input   io_sel_negative,
  input   io_sel_positive,
  input   io_sel_double_negative,
  input   io_sel_double_positive,
  input   io_x,
  input   io_x_sub,
  output  io_p
);
  wire  _io_p_T_2 = ~(io_sel_negative & ~io_x); // @[RS.scala 18:11]
  wire  _io_p_T_6 = _io_p_T_2 & ~(io_sel_double_negative & ~io_x_sub); // @[RS.scala 19:9]
  wire  _io_p_T_9 = _io_p_T_6 & ~(io_sel_positive & io_x); // @[RS.scala 20:9]
  wire  _io_p_T_12 = _io_p_T_9 & ~(io_sel_double_positive & io_x_sub); // @[RS.scala 21:9]
  assign io_p = ~_io_p_T_12; // @[RS.scala 18:9]
endmodule
module BOOTH_S(
  output       io_sel_negative,
  output       io_sel_positive,
  output       io_sel_double_negative,
  output       io_sel_double_positive,
  input  [2:0] io_src
);
  wire  y_add = io_src[2]; // @[BOOTH_S.scala 14:23]
  wire  y = io_src[1]; // @[BOOTH_S.scala 15:23]
  wire  y_sub = io_src[0]; // @[BOOTH_S.scala 16:23]
  wire  _io_sel_negative_T = ~y_sub; // @[BOOTH_S.scala 17:37]
  wire  _io_sel_negative_T_2 = ~y; // @[BOOTH_S.scala 17:46]
  wire  _io_sel_negative_T_4 = y & ~y_sub | ~y & y_sub; // @[BOOTH_S.scala 17:44]
  wire  _io_sel_positive_T = ~y_add; // @[BOOTH_S.scala 18:24]
  assign io_sel_negative = y_add & (y & ~y_sub | ~y & y_sub); // @[BOOTH_S.scala 17:30]
  assign io_sel_positive = ~y_add & _io_sel_negative_T_4; // @[BOOTH_S.scala 18:31]
  assign io_sel_double_negative = y_add & _io_sel_negative_T_2 & _io_sel_negative_T; // @[BOOTH_S.scala 19:42]
  assign io_sel_double_positive = _io_sel_positive_T & y & y_sub; // @[BOOTH_S.scala 20:42]
endmodule
module BOOTH_gen(
  input  [131:0] io_x,
  input  [2:0]   io_y,
  output [131:0] io_out
);
  wire  RS_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_1_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_1_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_1_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_1_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_1_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_1_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_1_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_2_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_2_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_2_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_2_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_2_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_2_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_2_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_3_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_3_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_3_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_3_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_3_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_3_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_3_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_4_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_4_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_4_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_4_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_4_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_4_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_4_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_5_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_5_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_5_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_5_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_5_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_5_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_5_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_6_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_6_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_6_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_6_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_6_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_6_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_6_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_7_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_7_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_7_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_7_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_7_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_7_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_7_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_8_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_8_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_8_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_8_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_8_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_8_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_8_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_9_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_9_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_9_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_9_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_9_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_9_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_9_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_10_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_10_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_10_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_10_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_10_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_10_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_10_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_11_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_11_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_11_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_11_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_11_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_11_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_11_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_12_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_12_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_12_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_12_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_12_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_12_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_12_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_13_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_13_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_13_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_13_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_13_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_13_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_13_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_14_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_14_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_14_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_14_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_14_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_14_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_14_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_15_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_15_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_15_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_15_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_15_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_15_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_15_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_16_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_16_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_16_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_16_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_16_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_16_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_16_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_17_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_17_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_17_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_17_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_17_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_17_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_17_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_18_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_18_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_18_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_18_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_18_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_18_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_18_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_19_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_19_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_19_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_19_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_19_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_19_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_19_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_20_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_20_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_20_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_20_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_20_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_20_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_20_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_21_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_21_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_21_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_21_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_21_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_21_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_21_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_22_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_22_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_22_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_22_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_22_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_22_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_22_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_23_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_23_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_23_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_23_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_23_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_23_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_23_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_24_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_24_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_24_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_24_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_24_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_24_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_24_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_25_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_25_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_25_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_25_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_25_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_25_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_25_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_26_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_26_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_26_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_26_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_26_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_26_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_26_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_27_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_27_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_27_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_27_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_27_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_27_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_27_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_28_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_28_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_28_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_28_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_28_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_28_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_28_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_29_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_29_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_29_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_29_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_29_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_29_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_29_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_30_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_30_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_30_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_30_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_30_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_30_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_30_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_31_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_31_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_31_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_31_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_31_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_31_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_31_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_32_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_32_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_32_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_32_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_32_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_32_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_32_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_33_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_33_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_33_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_33_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_33_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_33_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_33_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_34_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_34_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_34_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_34_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_34_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_34_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_34_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_35_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_35_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_35_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_35_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_35_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_35_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_35_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_36_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_36_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_36_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_36_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_36_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_36_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_36_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_37_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_37_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_37_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_37_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_37_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_37_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_37_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_38_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_38_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_38_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_38_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_38_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_38_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_38_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_39_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_39_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_39_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_39_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_39_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_39_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_39_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_40_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_40_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_40_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_40_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_40_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_40_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_40_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_41_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_41_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_41_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_41_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_41_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_41_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_41_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_42_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_42_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_42_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_42_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_42_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_42_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_42_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_43_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_43_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_43_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_43_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_43_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_43_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_43_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_44_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_44_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_44_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_44_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_44_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_44_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_44_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_45_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_45_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_45_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_45_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_45_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_45_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_45_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_46_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_46_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_46_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_46_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_46_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_46_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_46_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_47_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_47_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_47_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_47_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_47_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_47_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_47_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_48_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_48_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_48_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_48_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_48_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_48_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_48_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_49_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_49_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_49_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_49_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_49_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_49_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_49_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_50_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_50_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_50_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_50_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_50_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_50_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_50_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_51_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_51_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_51_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_51_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_51_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_51_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_51_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_52_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_52_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_52_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_52_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_52_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_52_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_52_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_53_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_53_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_53_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_53_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_53_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_53_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_53_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_54_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_54_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_54_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_54_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_54_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_54_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_54_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_55_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_55_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_55_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_55_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_55_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_55_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_55_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_56_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_56_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_56_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_56_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_56_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_56_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_56_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_57_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_57_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_57_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_57_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_57_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_57_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_57_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_58_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_58_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_58_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_58_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_58_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_58_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_58_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_59_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_59_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_59_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_59_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_59_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_59_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_59_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_60_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_60_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_60_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_60_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_60_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_60_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_60_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_61_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_61_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_61_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_61_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_61_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_61_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_61_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_62_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_62_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_62_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_62_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_62_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_62_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_62_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_63_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_63_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_63_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_63_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_63_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_63_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_63_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_64_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_64_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_64_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_64_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_64_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_64_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_64_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_65_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_65_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_65_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_65_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_65_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_65_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_65_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_66_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_66_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_66_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_66_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_66_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_66_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_66_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_67_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_67_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_67_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_67_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_67_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_67_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_67_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_68_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_68_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_68_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_68_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_68_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_68_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_68_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_69_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_69_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_69_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_69_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_69_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_69_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_69_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_70_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_70_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_70_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_70_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_70_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_70_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_70_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_71_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_71_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_71_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_71_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_71_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_71_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_71_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_72_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_72_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_72_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_72_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_72_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_72_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_72_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_73_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_73_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_73_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_73_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_73_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_73_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_73_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_74_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_74_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_74_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_74_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_74_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_74_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_74_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_75_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_75_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_75_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_75_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_75_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_75_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_75_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_76_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_76_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_76_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_76_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_76_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_76_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_76_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_77_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_77_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_77_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_77_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_77_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_77_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_77_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_78_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_78_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_78_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_78_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_78_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_78_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_78_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_79_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_79_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_79_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_79_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_79_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_79_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_79_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_80_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_80_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_80_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_80_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_80_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_80_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_80_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_81_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_81_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_81_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_81_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_81_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_81_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_81_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_82_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_82_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_82_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_82_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_82_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_82_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_82_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_83_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_83_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_83_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_83_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_83_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_83_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_83_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_84_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_84_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_84_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_84_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_84_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_84_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_84_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_85_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_85_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_85_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_85_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_85_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_85_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_85_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_86_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_86_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_86_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_86_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_86_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_86_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_86_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_87_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_87_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_87_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_87_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_87_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_87_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_87_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_88_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_88_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_88_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_88_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_88_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_88_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_88_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_89_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_89_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_89_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_89_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_89_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_89_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_89_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_90_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_90_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_90_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_90_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_90_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_90_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_90_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_91_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_91_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_91_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_91_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_91_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_91_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_91_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_92_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_92_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_92_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_92_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_92_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_92_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_92_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_93_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_93_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_93_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_93_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_93_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_93_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_93_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_94_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_94_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_94_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_94_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_94_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_94_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_94_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_95_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_95_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_95_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_95_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_95_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_95_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_95_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_96_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_96_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_96_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_96_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_96_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_96_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_96_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_97_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_97_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_97_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_97_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_97_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_97_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_97_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_98_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_98_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_98_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_98_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_98_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_98_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_98_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_99_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_99_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_99_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_99_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_99_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_99_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_99_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_100_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_100_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_100_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_100_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_100_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_100_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_100_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_101_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_101_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_101_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_101_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_101_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_101_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_101_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_102_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_102_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_102_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_102_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_102_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_102_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_102_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_103_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_103_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_103_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_103_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_103_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_103_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_103_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_104_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_104_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_104_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_104_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_104_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_104_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_104_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_105_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_105_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_105_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_105_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_105_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_105_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_105_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_106_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_106_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_106_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_106_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_106_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_106_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_106_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_107_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_107_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_107_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_107_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_107_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_107_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_107_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_108_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_108_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_108_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_108_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_108_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_108_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_108_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_109_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_109_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_109_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_109_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_109_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_109_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_109_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_110_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_110_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_110_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_110_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_110_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_110_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_110_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_111_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_111_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_111_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_111_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_111_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_111_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_111_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_112_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_112_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_112_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_112_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_112_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_112_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_112_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_113_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_113_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_113_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_113_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_113_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_113_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_113_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_114_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_114_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_114_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_114_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_114_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_114_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_114_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_115_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_115_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_115_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_115_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_115_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_115_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_115_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_116_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_116_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_116_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_116_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_116_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_116_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_116_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_117_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_117_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_117_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_117_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_117_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_117_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_117_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_118_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_118_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_118_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_118_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_118_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_118_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_118_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_119_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_119_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_119_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_119_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_119_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_119_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_119_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_120_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_120_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_120_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_120_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_120_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_120_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_120_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_121_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_121_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_121_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_121_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_121_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_121_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_121_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_122_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_122_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_122_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_122_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_122_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_122_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_122_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_123_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_123_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_123_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_123_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_123_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_123_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_123_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_124_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_124_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_124_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_124_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_124_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_124_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_124_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_125_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_125_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_125_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_125_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_125_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_125_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_125_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_126_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_126_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_126_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_126_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_126_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_126_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_126_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_127_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_127_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_127_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_127_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_127_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_127_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_127_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_128_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_128_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_128_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_128_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_128_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_128_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_128_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_129_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_129_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_129_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_129_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_129_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_129_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_129_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_130_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_130_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_130_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_130_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_130_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_130_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_130_io_p; // @[BOOTH_gen.scala 15:42]
  wire  RS_131_io_sel_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_131_io_sel_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_131_io_sel_double_negative; // @[BOOTH_gen.scala 15:42]
  wire  RS_131_io_sel_double_positive; // @[BOOTH_gen.scala 15:42]
  wire  RS_131_io_x; // @[BOOTH_gen.scala 15:42]
  wire  RS_131_io_x_sub; // @[BOOTH_gen.scala 15:42]
  wire  RS_131_io_p; // @[BOOTH_gen.scala 15:42]
  wire  BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:21]
  wire  BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:21]
  wire  BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:21]
  wire  BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:21]
  wire [2:0] BOOTH_S_io_src; // @[BOOTH_gen.scala 16:21]
  wire  r_1_p = RS_1_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_0_p = RS_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_3_p = RS_3_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_2_p = RS_2_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_5_p = RS_5_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_4_p = RS_4_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_7_p = RS_7_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_6_p = RS_6_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [7:0] io_out_lo_lo_lo_lo = {r_7_p,r_6_p,r_5_p,r_4_p,r_3_p,r_2_p,r_1_p,r_0_p}; // @[Cat.scala 31:58]
  wire  r_9_p = RS_9_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_8_p = RS_8_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_11_p = RS_11_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_10_p = RS_10_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_13_p = RS_13_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_12_p = RS_12_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_15_p = RS_15_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_14_p = RS_14_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_17_p = RS_17_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_16_p = RS_16_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_19_p = RS_19_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_18_p = RS_18_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_21_p = RS_21_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_20_p = RS_20_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_23_p = RS_23_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_22_p = RS_22_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [7:0] io_out_lo_lo_hi_lo = {r_23_p,r_22_p,r_21_p,r_20_p,r_19_p,r_18_p,r_17_p,r_16_p}; // @[Cat.scala 31:58]
  wire  r_25_p = RS_25_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_24_p = RS_24_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_27_p = RS_27_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_26_p = RS_26_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_29_p = RS_29_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_28_p = RS_28_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_32_p = RS_32_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_31_p = RS_31_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_30_p = RS_30_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [16:0] io_out_lo_lo_hi = {r_32_p,r_31_p,r_30_p,r_29_p,r_28_p,r_27_p,r_26_p,r_25_p,r_24_p,io_out_lo_lo_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] io_out_lo_lo = {io_out_lo_lo_hi,r_15_p,r_14_p,r_13_p,r_12_p,r_11_p,r_10_p,r_9_p,r_8_p,io_out_lo_lo_lo_lo}; // @[Cat.scala 31:58]
  wire  r_34_p = RS_34_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_33_p = RS_33_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_36_p = RS_36_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_35_p = RS_35_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_38_p = RS_38_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_37_p = RS_37_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_40_p = RS_40_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_39_p = RS_39_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [7:0] io_out_lo_hi_lo_lo = {r_40_p,r_39_p,r_38_p,r_37_p,r_36_p,r_35_p,r_34_p,r_33_p}; // @[Cat.scala 31:58]
  wire  r_42_p = RS_42_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_41_p = RS_41_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_44_p = RS_44_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_43_p = RS_43_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_46_p = RS_46_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_45_p = RS_45_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_48_p = RS_48_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_47_p = RS_47_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_50_p = RS_50_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_49_p = RS_49_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_52_p = RS_52_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_51_p = RS_51_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_54_p = RS_54_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_53_p = RS_53_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_56_p = RS_56_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_55_p = RS_55_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [7:0] io_out_lo_hi_hi_lo = {r_56_p,r_55_p,r_54_p,r_53_p,r_52_p,r_51_p,r_50_p,r_49_p}; // @[Cat.scala 31:58]
  wire  r_58_p = RS_58_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_57_p = RS_57_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_60_p = RS_60_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_59_p = RS_59_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_62_p = RS_62_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_61_p = RS_61_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_65_p = RS_65_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_64_p = RS_64_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_63_p = RS_63_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [16:0] io_out_lo_hi_hi = {r_65_p,r_64_p,r_63_p,r_62_p,r_61_p,r_60_p,r_59_p,r_58_p,r_57_p,io_out_lo_hi_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] io_out_lo_hi = {io_out_lo_hi_hi,r_48_p,r_47_p,r_46_p,r_45_p,r_44_p,r_43_p,r_42_p,r_41_p,io_out_lo_hi_lo_lo
    }; // @[Cat.scala 31:58]
  wire [65:0] io_out_lo = {io_out_lo_hi,io_out_lo_lo}; // @[Cat.scala 31:58]
  wire  r_67_p = RS_67_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_66_p = RS_66_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_69_p = RS_69_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_68_p = RS_68_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_71_p = RS_71_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_70_p = RS_70_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_73_p = RS_73_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_72_p = RS_72_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [7:0] io_out_hi_lo_lo_lo = {r_73_p,r_72_p,r_71_p,r_70_p,r_69_p,r_68_p,r_67_p,r_66_p}; // @[Cat.scala 31:58]
  wire  r_75_p = RS_75_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_74_p = RS_74_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_77_p = RS_77_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_76_p = RS_76_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_79_p = RS_79_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_78_p = RS_78_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_81_p = RS_81_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_80_p = RS_80_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_83_p = RS_83_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_82_p = RS_82_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_85_p = RS_85_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_84_p = RS_84_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_87_p = RS_87_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_86_p = RS_86_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_89_p = RS_89_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_88_p = RS_88_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [7:0] io_out_hi_lo_hi_lo = {r_89_p,r_88_p,r_87_p,r_86_p,r_85_p,r_84_p,r_83_p,r_82_p}; // @[Cat.scala 31:58]
  wire  r_91_p = RS_91_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_90_p = RS_90_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_93_p = RS_93_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_92_p = RS_92_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_95_p = RS_95_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_94_p = RS_94_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_98_p = RS_98_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_97_p = RS_97_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_96_p = RS_96_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [16:0] io_out_hi_lo_hi = {r_98_p,r_97_p,r_96_p,r_95_p,r_94_p,r_93_p,r_92_p,r_91_p,r_90_p,io_out_hi_lo_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] io_out_hi_lo = {io_out_hi_lo_hi,r_81_p,r_80_p,r_79_p,r_78_p,r_77_p,r_76_p,r_75_p,r_74_p,io_out_hi_lo_lo_lo
    }; // @[Cat.scala 31:58]
  wire  r_100_p = RS_100_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_99_p = RS_99_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_102_p = RS_102_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_101_p = RS_101_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_104_p = RS_104_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_103_p = RS_103_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_106_p = RS_106_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_105_p = RS_105_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [7:0] io_out_hi_hi_lo_lo = {r_106_p,r_105_p,r_104_p,r_103_p,r_102_p,r_101_p,r_100_p,r_99_p}; // @[Cat.scala 31:58]
  wire  r_108_p = RS_108_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_107_p = RS_107_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_110_p = RS_110_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_109_p = RS_109_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_112_p = RS_112_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_111_p = RS_111_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_114_p = RS_114_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_113_p = RS_113_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_116_p = RS_116_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_115_p = RS_115_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_118_p = RS_118_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_117_p = RS_117_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_120_p = RS_120_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_119_p = RS_119_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_122_p = RS_122_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_121_p = RS_121_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [7:0] io_out_hi_hi_hi_lo = {r_122_p,r_121_p,r_120_p,r_119_p,r_118_p,r_117_p,r_116_p,r_115_p}; // @[Cat.scala 31:58]
  wire  r_124_p = RS_124_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_123_p = RS_123_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_126_p = RS_126_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_125_p = RS_125_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_128_p = RS_128_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_127_p = RS_127_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_131_p = RS_131_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_130_p = RS_130_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire  r_129_p = RS_129_io_p; // @[BOOTH_gen.scala 15:{20,20}]
  wire [16:0] io_out_hi_hi_hi = {r_131_p,r_130_p,r_129_p,r_128_p,r_127_p,r_126_p,r_125_p,r_124_p,r_123_p,
    io_out_hi_hi_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] io_out_hi_hi = {io_out_hi_hi_hi,r_114_p,r_113_p,r_112_p,r_111_p,r_110_p,r_109_p,r_108_p,r_107_p,
    io_out_hi_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [65:0] io_out_hi = {io_out_hi_hi,io_out_hi_lo}; // @[Cat.scala 31:58]
  RS RS ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_io_sel_negative),
    .io_sel_positive(RS_io_sel_positive),
    .io_sel_double_negative(RS_io_sel_double_negative),
    .io_sel_double_positive(RS_io_sel_double_positive),
    .io_x(RS_io_x),
    .io_x_sub(RS_io_x_sub),
    .io_p(RS_io_p)
  );
  RS RS_1 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_1_io_sel_negative),
    .io_sel_positive(RS_1_io_sel_positive),
    .io_sel_double_negative(RS_1_io_sel_double_negative),
    .io_sel_double_positive(RS_1_io_sel_double_positive),
    .io_x(RS_1_io_x),
    .io_x_sub(RS_1_io_x_sub),
    .io_p(RS_1_io_p)
  );
  RS RS_2 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_2_io_sel_negative),
    .io_sel_positive(RS_2_io_sel_positive),
    .io_sel_double_negative(RS_2_io_sel_double_negative),
    .io_sel_double_positive(RS_2_io_sel_double_positive),
    .io_x(RS_2_io_x),
    .io_x_sub(RS_2_io_x_sub),
    .io_p(RS_2_io_p)
  );
  RS RS_3 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_3_io_sel_negative),
    .io_sel_positive(RS_3_io_sel_positive),
    .io_sel_double_negative(RS_3_io_sel_double_negative),
    .io_sel_double_positive(RS_3_io_sel_double_positive),
    .io_x(RS_3_io_x),
    .io_x_sub(RS_3_io_x_sub),
    .io_p(RS_3_io_p)
  );
  RS RS_4 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_4_io_sel_negative),
    .io_sel_positive(RS_4_io_sel_positive),
    .io_sel_double_negative(RS_4_io_sel_double_negative),
    .io_sel_double_positive(RS_4_io_sel_double_positive),
    .io_x(RS_4_io_x),
    .io_x_sub(RS_4_io_x_sub),
    .io_p(RS_4_io_p)
  );
  RS RS_5 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_5_io_sel_negative),
    .io_sel_positive(RS_5_io_sel_positive),
    .io_sel_double_negative(RS_5_io_sel_double_negative),
    .io_sel_double_positive(RS_5_io_sel_double_positive),
    .io_x(RS_5_io_x),
    .io_x_sub(RS_5_io_x_sub),
    .io_p(RS_5_io_p)
  );
  RS RS_6 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_6_io_sel_negative),
    .io_sel_positive(RS_6_io_sel_positive),
    .io_sel_double_negative(RS_6_io_sel_double_negative),
    .io_sel_double_positive(RS_6_io_sel_double_positive),
    .io_x(RS_6_io_x),
    .io_x_sub(RS_6_io_x_sub),
    .io_p(RS_6_io_p)
  );
  RS RS_7 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_7_io_sel_negative),
    .io_sel_positive(RS_7_io_sel_positive),
    .io_sel_double_negative(RS_7_io_sel_double_negative),
    .io_sel_double_positive(RS_7_io_sel_double_positive),
    .io_x(RS_7_io_x),
    .io_x_sub(RS_7_io_x_sub),
    .io_p(RS_7_io_p)
  );
  RS RS_8 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_8_io_sel_negative),
    .io_sel_positive(RS_8_io_sel_positive),
    .io_sel_double_negative(RS_8_io_sel_double_negative),
    .io_sel_double_positive(RS_8_io_sel_double_positive),
    .io_x(RS_8_io_x),
    .io_x_sub(RS_8_io_x_sub),
    .io_p(RS_8_io_p)
  );
  RS RS_9 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_9_io_sel_negative),
    .io_sel_positive(RS_9_io_sel_positive),
    .io_sel_double_negative(RS_9_io_sel_double_negative),
    .io_sel_double_positive(RS_9_io_sel_double_positive),
    .io_x(RS_9_io_x),
    .io_x_sub(RS_9_io_x_sub),
    .io_p(RS_9_io_p)
  );
  RS RS_10 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_10_io_sel_negative),
    .io_sel_positive(RS_10_io_sel_positive),
    .io_sel_double_negative(RS_10_io_sel_double_negative),
    .io_sel_double_positive(RS_10_io_sel_double_positive),
    .io_x(RS_10_io_x),
    .io_x_sub(RS_10_io_x_sub),
    .io_p(RS_10_io_p)
  );
  RS RS_11 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_11_io_sel_negative),
    .io_sel_positive(RS_11_io_sel_positive),
    .io_sel_double_negative(RS_11_io_sel_double_negative),
    .io_sel_double_positive(RS_11_io_sel_double_positive),
    .io_x(RS_11_io_x),
    .io_x_sub(RS_11_io_x_sub),
    .io_p(RS_11_io_p)
  );
  RS RS_12 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_12_io_sel_negative),
    .io_sel_positive(RS_12_io_sel_positive),
    .io_sel_double_negative(RS_12_io_sel_double_negative),
    .io_sel_double_positive(RS_12_io_sel_double_positive),
    .io_x(RS_12_io_x),
    .io_x_sub(RS_12_io_x_sub),
    .io_p(RS_12_io_p)
  );
  RS RS_13 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_13_io_sel_negative),
    .io_sel_positive(RS_13_io_sel_positive),
    .io_sel_double_negative(RS_13_io_sel_double_negative),
    .io_sel_double_positive(RS_13_io_sel_double_positive),
    .io_x(RS_13_io_x),
    .io_x_sub(RS_13_io_x_sub),
    .io_p(RS_13_io_p)
  );
  RS RS_14 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_14_io_sel_negative),
    .io_sel_positive(RS_14_io_sel_positive),
    .io_sel_double_negative(RS_14_io_sel_double_negative),
    .io_sel_double_positive(RS_14_io_sel_double_positive),
    .io_x(RS_14_io_x),
    .io_x_sub(RS_14_io_x_sub),
    .io_p(RS_14_io_p)
  );
  RS RS_15 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_15_io_sel_negative),
    .io_sel_positive(RS_15_io_sel_positive),
    .io_sel_double_negative(RS_15_io_sel_double_negative),
    .io_sel_double_positive(RS_15_io_sel_double_positive),
    .io_x(RS_15_io_x),
    .io_x_sub(RS_15_io_x_sub),
    .io_p(RS_15_io_p)
  );
  RS RS_16 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_16_io_sel_negative),
    .io_sel_positive(RS_16_io_sel_positive),
    .io_sel_double_negative(RS_16_io_sel_double_negative),
    .io_sel_double_positive(RS_16_io_sel_double_positive),
    .io_x(RS_16_io_x),
    .io_x_sub(RS_16_io_x_sub),
    .io_p(RS_16_io_p)
  );
  RS RS_17 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_17_io_sel_negative),
    .io_sel_positive(RS_17_io_sel_positive),
    .io_sel_double_negative(RS_17_io_sel_double_negative),
    .io_sel_double_positive(RS_17_io_sel_double_positive),
    .io_x(RS_17_io_x),
    .io_x_sub(RS_17_io_x_sub),
    .io_p(RS_17_io_p)
  );
  RS RS_18 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_18_io_sel_negative),
    .io_sel_positive(RS_18_io_sel_positive),
    .io_sel_double_negative(RS_18_io_sel_double_negative),
    .io_sel_double_positive(RS_18_io_sel_double_positive),
    .io_x(RS_18_io_x),
    .io_x_sub(RS_18_io_x_sub),
    .io_p(RS_18_io_p)
  );
  RS RS_19 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_19_io_sel_negative),
    .io_sel_positive(RS_19_io_sel_positive),
    .io_sel_double_negative(RS_19_io_sel_double_negative),
    .io_sel_double_positive(RS_19_io_sel_double_positive),
    .io_x(RS_19_io_x),
    .io_x_sub(RS_19_io_x_sub),
    .io_p(RS_19_io_p)
  );
  RS RS_20 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_20_io_sel_negative),
    .io_sel_positive(RS_20_io_sel_positive),
    .io_sel_double_negative(RS_20_io_sel_double_negative),
    .io_sel_double_positive(RS_20_io_sel_double_positive),
    .io_x(RS_20_io_x),
    .io_x_sub(RS_20_io_x_sub),
    .io_p(RS_20_io_p)
  );
  RS RS_21 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_21_io_sel_negative),
    .io_sel_positive(RS_21_io_sel_positive),
    .io_sel_double_negative(RS_21_io_sel_double_negative),
    .io_sel_double_positive(RS_21_io_sel_double_positive),
    .io_x(RS_21_io_x),
    .io_x_sub(RS_21_io_x_sub),
    .io_p(RS_21_io_p)
  );
  RS RS_22 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_22_io_sel_negative),
    .io_sel_positive(RS_22_io_sel_positive),
    .io_sel_double_negative(RS_22_io_sel_double_negative),
    .io_sel_double_positive(RS_22_io_sel_double_positive),
    .io_x(RS_22_io_x),
    .io_x_sub(RS_22_io_x_sub),
    .io_p(RS_22_io_p)
  );
  RS RS_23 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_23_io_sel_negative),
    .io_sel_positive(RS_23_io_sel_positive),
    .io_sel_double_negative(RS_23_io_sel_double_negative),
    .io_sel_double_positive(RS_23_io_sel_double_positive),
    .io_x(RS_23_io_x),
    .io_x_sub(RS_23_io_x_sub),
    .io_p(RS_23_io_p)
  );
  RS RS_24 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_24_io_sel_negative),
    .io_sel_positive(RS_24_io_sel_positive),
    .io_sel_double_negative(RS_24_io_sel_double_negative),
    .io_sel_double_positive(RS_24_io_sel_double_positive),
    .io_x(RS_24_io_x),
    .io_x_sub(RS_24_io_x_sub),
    .io_p(RS_24_io_p)
  );
  RS RS_25 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_25_io_sel_negative),
    .io_sel_positive(RS_25_io_sel_positive),
    .io_sel_double_negative(RS_25_io_sel_double_negative),
    .io_sel_double_positive(RS_25_io_sel_double_positive),
    .io_x(RS_25_io_x),
    .io_x_sub(RS_25_io_x_sub),
    .io_p(RS_25_io_p)
  );
  RS RS_26 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_26_io_sel_negative),
    .io_sel_positive(RS_26_io_sel_positive),
    .io_sel_double_negative(RS_26_io_sel_double_negative),
    .io_sel_double_positive(RS_26_io_sel_double_positive),
    .io_x(RS_26_io_x),
    .io_x_sub(RS_26_io_x_sub),
    .io_p(RS_26_io_p)
  );
  RS RS_27 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_27_io_sel_negative),
    .io_sel_positive(RS_27_io_sel_positive),
    .io_sel_double_negative(RS_27_io_sel_double_negative),
    .io_sel_double_positive(RS_27_io_sel_double_positive),
    .io_x(RS_27_io_x),
    .io_x_sub(RS_27_io_x_sub),
    .io_p(RS_27_io_p)
  );
  RS RS_28 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_28_io_sel_negative),
    .io_sel_positive(RS_28_io_sel_positive),
    .io_sel_double_negative(RS_28_io_sel_double_negative),
    .io_sel_double_positive(RS_28_io_sel_double_positive),
    .io_x(RS_28_io_x),
    .io_x_sub(RS_28_io_x_sub),
    .io_p(RS_28_io_p)
  );
  RS RS_29 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_29_io_sel_negative),
    .io_sel_positive(RS_29_io_sel_positive),
    .io_sel_double_negative(RS_29_io_sel_double_negative),
    .io_sel_double_positive(RS_29_io_sel_double_positive),
    .io_x(RS_29_io_x),
    .io_x_sub(RS_29_io_x_sub),
    .io_p(RS_29_io_p)
  );
  RS RS_30 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_30_io_sel_negative),
    .io_sel_positive(RS_30_io_sel_positive),
    .io_sel_double_negative(RS_30_io_sel_double_negative),
    .io_sel_double_positive(RS_30_io_sel_double_positive),
    .io_x(RS_30_io_x),
    .io_x_sub(RS_30_io_x_sub),
    .io_p(RS_30_io_p)
  );
  RS RS_31 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_31_io_sel_negative),
    .io_sel_positive(RS_31_io_sel_positive),
    .io_sel_double_negative(RS_31_io_sel_double_negative),
    .io_sel_double_positive(RS_31_io_sel_double_positive),
    .io_x(RS_31_io_x),
    .io_x_sub(RS_31_io_x_sub),
    .io_p(RS_31_io_p)
  );
  RS RS_32 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_32_io_sel_negative),
    .io_sel_positive(RS_32_io_sel_positive),
    .io_sel_double_negative(RS_32_io_sel_double_negative),
    .io_sel_double_positive(RS_32_io_sel_double_positive),
    .io_x(RS_32_io_x),
    .io_x_sub(RS_32_io_x_sub),
    .io_p(RS_32_io_p)
  );
  RS RS_33 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_33_io_sel_negative),
    .io_sel_positive(RS_33_io_sel_positive),
    .io_sel_double_negative(RS_33_io_sel_double_negative),
    .io_sel_double_positive(RS_33_io_sel_double_positive),
    .io_x(RS_33_io_x),
    .io_x_sub(RS_33_io_x_sub),
    .io_p(RS_33_io_p)
  );
  RS RS_34 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_34_io_sel_negative),
    .io_sel_positive(RS_34_io_sel_positive),
    .io_sel_double_negative(RS_34_io_sel_double_negative),
    .io_sel_double_positive(RS_34_io_sel_double_positive),
    .io_x(RS_34_io_x),
    .io_x_sub(RS_34_io_x_sub),
    .io_p(RS_34_io_p)
  );
  RS RS_35 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_35_io_sel_negative),
    .io_sel_positive(RS_35_io_sel_positive),
    .io_sel_double_negative(RS_35_io_sel_double_negative),
    .io_sel_double_positive(RS_35_io_sel_double_positive),
    .io_x(RS_35_io_x),
    .io_x_sub(RS_35_io_x_sub),
    .io_p(RS_35_io_p)
  );
  RS RS_36 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_36_io_sel_negative),
    .io_sel_positive(RS_36_io_sel_positive),
    .io_sel_double_negative(RS_36_io_sel_double_negative),
    .io_sel_double_positive(RS_36_io_sel_double_positive),
    .io_x(RS_36_io_x),
    .io_x_sub(RS_36_io_x_sub),
    .io_p(RS_36_io_p)
  );
  RS RS_37 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_37_io_sel_negative),
    .io_sel_positive(RS_37_io_sel_positive),
    .io_sel_double_negative(RS_37_io_sel_double_negative),
    .io_sel_double_positive(RS_37_io_sel_double_positive),
    .io_x(RS_37_io_x),
    .io_x_sub(RS_37_io_x_sub),
    .io_p(RS_37_io_p)
  );
  RS RS_38 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_38_io_sel_negative),
    .io_sel_positive(RS_38_io_sel_positive),
    .io_sel_double_negative(RS_38_io_sel_double_negative),
    .io_sel_double_positive(RS_38_io_sel_double_positive),
    .io_x(RS_38_io_x),
    .io_x_sub(RS_38_io_x_sub),
    .io_p(RS_38_io_p)
  );
  RS RS_39 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_39_io_sel_negative),
    .io_sel_positive(RS_39_io_sel_positive),
    .io_sel_double_negative(RS_39_io_sel_double_negative),
    .io_sel_double_positive(RS_39_io_sel_double_positive),
    .io_x(RS_39_io_x),
    .io_x_sub(RS_39_io_x_sub),
    .io_p(RS_39_io_p)
  );
  RS RS_40 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_40_io_sel_negative),
    .io_sel_positive(RS_40_io_sel_positive),
    .io_sel_double_negative(RS_40_io_sel_double_negative),
    .io_sel_double_positive(RS_40_io_sel_double_positive),
    .io_x(RS_40_io_x),
    .io_x_sub(RS_40_io_x_sub),
    .io_p(RS_40_io_p)
  );
  RS RS_41 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_41_io_sel_negative),
    .io_sel_positive(RS_41_io_sel_positive),
    .io_sel_double_negative(RS_41_io_sel_double_negative),
    .io_sel_double_positive(RS_41_io_sel_double_positive),
    .io_x(RS_41_io_x),
    .io_x_sub(RS_41_io_x_sub),
    .io_p(RS_41_io_p)
  );
  RS RS_42 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_42_io_sel_negative),
    .io_sel_positive(RS_42_io_sel_positive),
    .io_sel_double_negative(RS_42_io_sel_double_negative),
    .io_sel_double_positive(RS_42_io_sel_double_positive),
    .io_x(RS_42_io_x),
    .io_x_sub(RS_42_io_x_sub),
    .io_p(RS_42_io_p)
  );
  RS RS_43 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_43_io_sel_negative),
    .io_sel_positive(RS_43_io_sel_positive),
    .io_sel_double_negative(RS_43_io_sel_double_negative),
    .io_sel_double_positive(RS_43_io_sel_double_positive),
    .io_x(RS_43_io_x),
    .io_x_sub(RS_43_io_x_sub),
    .io_p(RS_43_io_p)
  );
  RS RS_44 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_44_io_sel_negative),
    .io_sel_positive(RS_44_io_sel_positive),
    .io_sel_double_negative(RS_44_io_sel_double_negative),
    .io_sel_double_positive(RS_44_io_sel_double_positive),
    .io_x(RS_44_io_x),
    .io_x_sub(RS_44_io_x_sub),
    .io_p(RS_44_io_p)
  );
  RS RS_45 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_45_io_sel_negative),
    .io_sel_positive(RS_45_io_sel_positive),
    .io_sel_double_negative(RS_45_io_sel_double_negative),
    .io_sel_double_positive(RS_45_io_sel_double_positive),
    .io_x(RS_45_io_x),
    .io_x_sub(RS_45_io_x_sub),
    .io_p(RS_45_io_p)
  );
  RS RS_46 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_46_io_sel_negative),
    .io_sel_positive(RS_46_io_sel_positive),
    .io_sel_double_negative(RS_46_io_sel_double_negative),
    .io_sel_double_positive(RS_46_io_sel_double_positive),
    .io_x(RS_46_io_x),
    .io_x_sub(RS_46_io_x_sub),
    .io_p(RS_46_io_p)
  );
  RS RS_47 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_47_io_sel_negative),
    .io_sel_positive(RS_47_io_sel_positive),
    .io_sel_double_negative(RS_47_io_sel_double_negative),
    .io_sel_double_positive(RS_47_io_sel_double_positive),
    .io_x(RS_47_io_x),
    .io_x_sub(RS_47_io_x_sub),
    .io_p(RS_47_io_p)
  );
  RS RS_48 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_48_io_sel_negative),
    .io_sel_positive(RS_48_io_sel_positive),
    .io_sel_double_negative(RS_48_io_sel_double_negative),
    .io_sel_double_positive(RS_48_io_sel_double_positive),
    .io_x(RS_48_io_x),
    .io_x_sub(RS_48_io_x_sub),
    .io_p(RS_48_io_p)
  );
  RS RS_49 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_49_io_sel_negative),
    .io_sel_positive(RS_49_io_sel_positive),
    .io_sel_double_negative(RS_49_io_sel_double_negative),
    .io_sel_double_positive(RS_49_io_sel_double_positive),
    .io_x(RS_49_io_x),
    .io_x_sub(RS_49_io_x_sub),
    .io_p(RS_49_io_p)
  );
  RS RS_50 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_50_io_sel_negative),
    .io_sel_positive(RS_50_io_sel_positive),
    .io_sel_double_negative(RS_50_io_sel_double_negative),
    .io_sel_double_positive(RS_50_io_sel_double_positive),
    .io_x(RS_50_io_x),
    .io_x_sub(RS_50_io_x_sub),
    .io_p(RS_50_io_p)
  );
  RS RS_51 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_51_io_sel_negative),
    .io_sel_positive(RS_51_io_sel_positive),
    .io_sel_double_negative(RS_51_io_sel_double_negative),
    .io_sel_double_positive(RS_51_io_sel_double_positive),
    .io_x(RS_51_io_x),
    .io_x_sub(RS_51_io_x_sub),
    .io_p(RS_51_io_p)
  );
  RS RS_52 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_52_io_sel_negative),
    .io_sel_positive(RS_52_io_sel_positive),
    .io_sel_double_negative(RS_52_io_sel_double_negative),
    .io_sel_double_positive(RS_52_io_sel_double_positive),
    .io_x(RS_52_io_x),
    .io_x_sub(RS_52_io_x_sub),
    .io_p(RS_52_io_p)
  );
  RS RS_53 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_53_io_sel_negative),
    .io_sel_positive(RS_53_io_sel_positive),
    .io_sel_double_negative(RS_53_io_sel_double_negative),
    .io_sel_double_positive(RS_53_io_sel_double_positive),
    .io_x(RS_53_io_x),
    .io_x_sub(RS_53_io_x_sub),
    .io_p(RS_53_io_p)
  );
  RS RS_54 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_54_io_sel_negative),
    .io_sel_positive(RS_54_io_sel_positive),
    .io_sel_double_negative(RS_54_io_sel_double_negative),
    .io_sel_double_positive(RS_54_io_sel_double_positive),
    .io_x(RS_54_io_x),
    .io_x_sub(RS_54_io_x_sub),
    .io_p(RS_54_io_p)
  );
  RS RS_55 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_55_io_sel_negative),
    .io_sel_positive(RS_55_io_sel_positive),
    .io_sel_double_negative(RS_55_io_sel_double_negative),
    .io_sel_double_positive(RS_55_io_sel_double_positive),
    .io_x(RS_55_io_x),
    .io_x_sub(RS_55_io_x_sub),
    .io_p(RS_55_io_p)
  );
  RS RS_56 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_56_io_sel_negative),
    .io_sel_positive(RS_56_io_sel_positive),
    .io_sel_double_negative(RS_56_io_sel_double_negative),
    .io_sel_double_positive(RS_56_io_sel_double_positive),
    .io_x(RS_56_io_x),
    .io_x_sub(RS_56_io_x_sub),
    .io_p(RS_56_io_p)
  );
  RS RS_57 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_57_io_sel_negative),
    .io_sel_positive(RS_57_io_sel_positive),
    .io_sel_double_negative(RS_57_io_sel_double_negative),
    .io_sel_double_positive(RS_57_io_sel_double_positive),
    .io_x(RS_57_io_x),
    .io_x_sub(RS_57_io_x_sub),
    .io_p(RS_57_io_p)
  );
  RS RS_58 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_58_io_sel_negative),
    .io_sel_positive(RS_58_io_sel_positive),
    .io_sel_double_negative(RS_58_io_sel_double_negative),
    .io_sel_double_positive(RS_58_io_sel_double_positive),
    .io_x(RS_58_io_x),
    .io_x_sub(RS_58_io_x_sub),
    .io_p(RS_58_io_p)
  );
  RS RS_59 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_59_io_sel_negative),
    .io_sel_positive(RS_59_io_sel_positive),
    .io_sel_double_negative(RS_59_io_sel_double_negative),
    .io_sel_double_positive(RS_59_io_sel_double_positive),
    .io_x(RS_59_io_x),
    .io_x_sub(RS_59_io_x_sub),
    .io_p(RS_59_io_p)
  );
  RS RS_60 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_60_io_sel_negative),
    .io_sel_positive(RS_60_io_sel_positive),
    .io_sel_double_negative(RS_60_io_sel_double_negative),
    .io_sel_double_positive(RS_60_io_sel_double_positive),
    .io_x(RS_60_io_x),
    .io_x_sub(RS_60_io_x_sub),
    .io_p(RS_60_io_p)
  );
  RS RS_61 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_61_io_sel_negative),
    .io_sel_positive(RS_61_io_sel_positive),
    .io_sel_double_negative(RS_61_io_sel_double_negative),
    .io_sel_double_positive(RS_61_io_sel_double_positive),
    .io_x(RS_61_io_x),
    .io_x_sub(RS_61_io_x_sub),
    .io_p(RS_61_io_p)
  );
  RS RS_62 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_62_io_sel_negative),
    .io_sel_positive(RS_62_io_sel_positive),
    .io_sel_double_negative(RS_62_io_sel_double_negative),
    .io_sel_double_positive(RS_62_io_sel_double_positive),
    .io_x(RS_62_io_x),
    .io_x_sub(RS_62_io_x_sub),
    .io_p(RS_62_io_p)
  );
  RS RS_63 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_63_io_sel_negative),
    .io_sel_positive(RS_63_io_sel_positive),
    .io_sel_double_negative(RS_63_io_sel_double_negative),
    .io_sel_double_positive(RS_63_io_sel_double_positive),
    .io_x(RS_63_io_x),
    .io_x_sub(RS_63_io_x_sub),
    .io_p(RS_63_io_p)
  );
  RS RS_64 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_64_io_sel_negative),
    .io_sel_positive(RS_64_io_sel_positive),
    .io_sel_double_negative(RS_64_io_sel_double_negative),
    .io_sel_double_positive(RS_64_io_sel_double_positive),
    .io_x(RS_64_io_x),
    .io_x_sub(RS_64_io_x_sub),
    .io_p(RS_64_io_p)
  );
  RS RS_65 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_65_io_sel_negative),
    .io_sel_positive(RS_65_io_sel_positive),
    .io_sel_double_negative(RS_65_io_sel_double_negative),
    .io_sel_double_positive(RS_65_io_sel_double_positive),
    .io_x(RS_65_io_x),
    .io_x_sub(RS_65_io_x_sub),
    .io_p(RS_65_io_p)
  );
  RS RS_66 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_66_io_sel_negative),
    .io_sel_positive(RS_66_io_sel_positive),
    .io_sel_double_negative(RS_66_io_sel_double_negative),
    .io_sel_double_positive(RS_66_io_sel_double_positive),
    .io_x(RS_66_io_x),
    .io_x_sub(RS_66_io_x_sub),
    .io_p(RS_66_io_p)
  );
  RS RS_67 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_67_io_sel_negative),
    .io_sel_positive(RS_67_io_sel_positive),
    .io_sel_double_negative(RS_67_io_sel_double_negative),
    .io_sel_double_positive(RS_67_io_sel_double_positive),
    .io_x(RS_67_io_x),
    .io_x_sub(RS_67_io_x_sub),
    .io_p(RS_67_io_p)
  );
  RS RS_68 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_68_io_sel_negative),
    .io_sel_positive(RS_68_io_sel_positive),
    .io_sel_double_negative(RS_68_io_sel_double_negative),
    .io_sel_double_positive(RS_68_io_sel_double_positive),
    .io_x(RS_68_io_x),
    .io_x_sub(RS_68_io_x_sub),
    .io_p(RS_68_io_p)
  );
  RS RS_69 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_69_io_sel_negative),
    .io_sel_positive(RS_69_io_sel_positive),
    .io_sel_double_negative(RS_69_io_sel_double_negative),
    .io_sel_double_positive(RS_69_io_sel_double_positive),
    .io_x(RS_69_io_x),
    .io_x_sub(RS_69_io_x_sub),
    .io_p(RS_69_io_p)
  );
  RS RS_70 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_70_io_sel_negative),
    .io_sel_positive(RS_70_io_sel_positive),
    .io_sel_double_negative(RS_70_io_sel_double_negative),
    .io_sel_double_positive(RS_70_io_sel_double_positive),
    .io_x(RS_70_io_x),
    .io_x_sub(RS_70_io_x_sub),
    .io_p(RS_70_io_p)
  );
  RS RS_71 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_71_io_sel_negative),
    .io_sel_positive(RS_71_io_sel_positive),
    .io_sel_double_negative(RS_71_io_sel_double_negative),
    .io_sel_double_positive(RS_71_io_sel_double_positive),
    .io_x(RS_71_io_x),
    .io_x_sub(RS_71_io_x_sub),
    .io_p(RS_71_io_p)
  );
  RS RS_72 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_72_io_sel_negative),
    .io_sel_positive(RS_72_io_sel_positive),
    .io_sel_double_negative(RS_72_io_sel_double_negative),
    .io_sel_double_positive(RS_72_io_sel_double_positive),
    .io_x(RS_72_io_x),
    .io_x_sub(RS_72_io_x_sub),
    .io_p(RS_72_io_p)
  );
  RS RS_73 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_73_io_sel_negative),
    .io_sel_positive(RS_73_io_sel_positive),
    .io_sel_double_negative(RS_73_io_sel_double_negative),
    .io_sel_double_positive(RS_73_io_sel_double_positive),
    .io_x(RS_73_io_x),
    .io_x_sub(RS_73_io_x_sub),
    .io_p(RS_73_io_p)
  );
  RS RS_74 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_74_io_sel_negative),
    .io_sel_positive(RS_74_io_sel_positive),
    .io_sel_double_negative(RS_74_io_sel_double_negative),
    .io_sel_double_positive(RS_74_io_sel_double_positive),
    .io_x(RS_74_io_x),
    .io_x_sub(RS_74_io_x_sub),
    .io_p(RS_74_io_p)
  );
  RS RS_75 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_75_io_sel_negative),
    .io_sel_positive(RS_75_io_sel_positive),
    .io_sel_double_negative(RS_75_io_sel_double_negative),
    .io_sel_double_positive(RS_75_io_sel_double_positive),
    .io_x(RS_75_io_x),
    .io_x_sub(RS_75_io_x_sub),
    .io_p(RS_75_io_p)
  );
  RS RS_76 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_76_io_sel_negative),
    .io_sel_positive(RS_76_io_sel_positive),
    .io_sel_double_negative(RS_76_io_sel_double_negative),
    .io_sel_double_positive(RS_76_io_sel_double_positive),
    .io_x(RS_76_io_x),
    .io_x_sub(RS_76_io_x_sub),
    .io_p(RS_76_io_p)
  );
  RS RS_77 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_77_io_sel_negative),
    .io_sel_positive(RS_77_io_sel_positive),
    .io_sel_double_negative(RS_77_io_sel_double_negative),
    .io_sel_double_positive(RS_77_io_sel_double_positive),
    .io_x(RS_77_io_x),
    .io_x_sub(RS_77_io_x_sub),
    .io_p(RS_77_io_p)
  );
  RS RS_78 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_78_io_sel_negative),
    .io_sel_positive(RS_78_io_sel_positive),
    .io_sel_double_negative(RS_78_io_sel_double_negative),
    .io_sel_double_positive(RS_78_io_sel_double_positive),
    .io_x(RS_78_io_x),
    .io_x_sub(RS_78_io_x_sub),
    .io_p(RS_78_io_p)
  );
  RS RS_79 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_79_io_sel_negative),
    .io_sel_positive(RS_79_io_sel_positive),
    .io_sel_double_negative(RS_79_io_sel_double_negative),
    .io_sel_double_positive(RS_79_io_sel_double_positive),
    .io_x(RS_79_io_x),
    .io_x_sub(RS_79_io_x_sub),
    .io_p(RS_79_io_p)
  );
  RS RS_80 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_80_io_sel_negative),
    .io_sel_positive(RS_80_io_sel_positive),
    .io_sel_double_negative(RS_80_io_sel_double_negative),
    .io_sel_double_positive(RS_80_io_sel_double_positive),
    .io_x(RS_80_io_x),
    .io_x_sub(RS_80_io_x_sub),
    .io_p(RS_80_io_p)
  );
  RS RS_81 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_81_io_sel_negative),
    .io_sel_positive(RS_81_io_sel_positive),
    .io_sel_double_negative(RS_81_io_sel_double_negative),
    .io_sel_double_positive(RS_81_io_sel_double_positive),
    .io_x(RS_81_io_x),
    .io_x_sub(RS_81_io_x_sub),
    .io_p(RS_81_io_p)
  );
  RS RS_82 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_82_io_sel_negative),
    .io_sel_positive(RS_82_io_sel_positive),
    .io_sel_double_negative(RS_82_io_sel_double_negative),
    .io_sel_double_positive(RS_82_io_sel_double_positive),
    .io_x(RS_82_io_x),
    .io_x_sub(RS_82_io_x_sub),
    .io_p(RS_82_io_p)
  );
  RS RS_83 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_83_io_sel_negative),
    .io_sel_positive(RS_83_io_sel_positive),
    .io_sel_double_negative(RS_83_io_sel_double_negative),
    .io_sel_double_positive(RS_83_io_sel_double_positive),
    .io_x(RS_83_io_x),
    .io_x_sub(RS_83_io_x_sub),
    .io_p(RS_83_io_p)
  );
  RS RS_84 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_84_io_sel_negative),
    .io_sel_positive(RS_84_io_sel_positive),
    .io_sel_double_negative(RS_84_io_sel_double_negative),
    .io_sel_double_positive(RS_84_io_sel_double_positive),
    .io_x(RS_84_io_x),
    .io_x_sub(RS_84_io_x_sub),
    .io_p(RS_84_io_p)
  );
  RS RS_85 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_85_io_sel_negative),
    .io_sel_positive(RS_85_io_sel_positive),
    .io_sel_double_negative(RS_85_io_sel_double_negative),
    .io_sel_double_positive(RS_85_io_sel_double_positive),
    .io_x(RS_85_io_x),
    .io_x_sub(RS_85_io_x_sub),
    .io_p(RS_85_io_p)
  );
  RS RS_86 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_86_io_sel_negative),
    .io_sel_positive(RS_86_io_sel_positive),
    .io_sel_double_negative(RS_86_io_sel_double_negative),
    .io_sel_double_positive(RS_86_io_sel_double_positive),
    .io_x(RS_86_io_x),
    .io_x_sub(RS_86_io_x_sub),
    .io_p(RS_86_io_p)
  );
  RS RS_87 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_87_io_sel_negative),
    .io_sel_positive(RS_87_io_sel_positive),
    .io_sel_double_negative(RS_87_io_sel_double_negative),
    .io_sel_double_positive(RS_87_io_sel_double_positive),
    .io_x(RS_87_io_x),
    .io_x_sub(RS_87_io_x_sub),
    .io_p(RS_87_io_p)
  );
  RS RS_88 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_88_io_sel_negative),
    .io_sel_positive(RS_88_io_sel_positive),
    .io_sel_double_negative(RS_88_io_sel_double_negative),
    .io_sel_double_positive(RS_88_io_sel_double_positive),
    .io_x(RS_88_io_x),
    .io_x_sub(RS_88_io_x_sub),
    .io_p(RS_88_io_p)
  );
  RS RS_89 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_89_io_sel_negative),
    .io_sel_positive(RS_89_io_sel_positive),
    .io_sel_double_negative(RS_89_io_sel_double_negative),
    .io_sel_double_positive(RS_89_io_sel_double_positive),
    .io_x(RS_89_io_x),
    .io_x_sub(RS_89_io_x_sub),
    .io_p(RS_89_io_p)
  );
  RS RS_90 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_90_io_sel_negative),
    .io_sel_positive(RS_90_io_sel_positive),
    .io_sel_double_negative(RS_90_io_sel_double_negative),
    .io_sel_double_positive(RS_90_io_sel_double_positive),
    .io_x(RS_90_io_x),
    .io_x_sub(RS_90_io_x_sub),
    .io_p(RS_90_io_p)
  );
  RS RS_91 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_91_io_sel_negative),
    .io_sel_positive(RS_91_io_sel_positive),
    .io_sel_double_negative(RS_91_io_sel_double_negative),
    .io_sel_double_positive(RS_91_io_sel_double_positive),
    .io_x(RS_91_io_x),
    .io_x_sub(RS_91_io_x_sub),
    .io_p(RS_91_io_p)
  );
  RS RS_92 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_92_io_sel_negative),
    .io_sel_positive(RS_92_io_sel_positive),
    .io_sel_double_negative(RS_92_io_sel_double_negative),
    .io_sel_double_positive(RS_92_io_sel_double_positive),
    .io_x(RS_92_io_x),
    .io_x_sub(RS_92_io_x_sub),
    .io_p(RS_92_io_p)
  );
  RS RS_93 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_93_io_sel_negative),
    .io_sel_positive(RS_93_io_sel_positive),
    .io_sel_double_negative(RS_93_io_sel_double_negative),
    .io_sel_double_positive(RS_93_io_sel_double_positive),
    .io_x(RS_93_io_x),
    .io_x_sub(RS_93_io_x_sub),
    .io_p(RS_93_io_p)
  );
  RS RS_94 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_94_io_sel_negative),
    .io_sel_positive(RS_94_io_sel_positive),
    .io_sel_double_negative(RS_94_io_sel_double_negative),
    .io_sel_double_positive(RS_94_io_sel_double_positive),
    .io_x(RS_94_io_x),
    .io_x_sub(RS_94_io_x_sub),
    .io_p(RS_94_io_p)
  );
  RS RS_95 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_95_io_sel_negative),
    .io_sel_positive(RS_95_io_sel_positive),
    .io_sel_double_negative(RS_95_io_sel_double_negative),
    .io_sel_double_positive(RS_95_io_sel_double_positive),
    .io_x(RS_95_io_x),
    .io_x_sub(RS_95_io_x_sub),
    .io_p(RS_95_io_p)
  );
  RS RS_96 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_96_io_sel_negative),
    .io_sel_positive(RS_96_io_sel_positive),
    .io_sel_double_negative(RS_96_io_sel_double_negative),
    .io_sel_double_positive(RS_96_io_sel_double_positive),
    .io_x(RS_96_io_x),
    .io_x_sub(RS_96_io_x_sub),
    .io_p(RS_96_io_p)
  );
  RS RS_97 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_97_io_sel_negative),
    .io_sel_positive(RS_97_io_sel_positive),
    .io_sel_double_negative(RS_97_io_sel_double_negative),
    .io_sel_double_positive(RS_97_io_sel_double_positive),
    .io_x(RS_97_io_x),
    .io_x_sub(RS_97_io_x_sub),
    .io_p(RS_97_io_p)
  );
  RS RS_98 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_98_io_sel_negative),
    .io_sel_positive(RS_98_io_sel_positive),
    .io_sel_double_negative(RS_98_io_sel_double_negative),
    .io_sel_double_positive(RS_98_io_sel_double_positive),
    .io_x(RS_98_io_x),
    .io_x_sub(RS_98_io_x_sub),
    .io_p(RS_98_io_p)
  );
  RS RS_99 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_99_io_sel_negative),
    .io_sel_positive(RS_99_io_sel_positive),
    .io_sel_double_negative(RS_99_io_sel_double_negative),
    .io_sel_double_positive(RS_99_io_sel_double_positive),
    .io_x(RS_99_io_x),
    .io_x_sub(RS_99_io_x_sub),
    .io_p(RS_99_io_p)
  );
  RS RS_100 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_100_io_sel_negative),
    .io_sel_positive(RS_100_io_sel_positive),
    .io_sel_double_negative(RS_100_io_sel_double_negative),
    .io_sel_double_positive(RS_100_io_sel_double_positive),
    .io_x(RS_100_io_x),
    .io_x_sub(RS_100_io_x_sub),
    .io_p(RS_100_io_p)
  );
  RS RS_101 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_101_io_sel_negative),
    .io_sel_positive(RS_101_io_sel_positive),
    .io_sel_double_negative(RS_101_io_sel_double_negative),
    .io_sel_double_positive(RS_101_io_sel_double_positive),
    .io_x(RS_101_io_x),
    .io_x_sub(RS_101_io_x_sub),
    .io_p(RS_101_io_p)
  );
  RS RS_102 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_102_io_sel_negative),
    .io_sel_positive(RS_102_io_sel_positive),
    .io_sel_double_negative(RS_102_io_sel_double_negative),
    .io_sel_double_positive(RS_102_io_sel_double_positive),
    .io_x(RS_102_io_x),
    .io_x_sub(RS_102_io_x_sub),
    .io_p(RS_102_io_p)
  );
  RS RS_103 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_103_io_sel_negative),
    .io_sel_positive(RS_103_io_sel_positive),
    .io_sel_double_negative(RS_103_io_sel_double_negative),
    .io_sel_double_positive(RS_103_io_sel_double_positive),
    .io_x(RS_103_io_x),
    .io_x_sub(RS_103_io_x_sub),
    .io_p(RS_103_io_p)
  );
  RS RS_104 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_104_io_sel_negative),
    .io_sel_positive(RS_104_io_sel_positive),
    .io_sel_double_negative(RS_104_io_sel_double_negative),
    .io_sel_double_positive(RS_104_io_sel_double_positive),
    .io_x(RS_104_io_x),
    .io_x_sub(RS_104_io_x_sub),
    .io_p(RS_104_io_p)
  );
  RS RS_105 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_105_io_sel_negative),
    .io_sel_positive(RS_105_io_sel_positive),
    .io_sel_double_negative(RS_105_io_sel_double_negative),
    .io_sel_double_positive(RS_105_io_sel_double_positive),
    .io_x(RS_105_io_x),
    .io_x_sub(RS_105_io_x_sub),
    .io_p(RS_105_io_p)
  );
  RS RS_106 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_106_io_sel_negative),
    .io_sel_positive(RS_106_io_sel_positive),
    .io_sel_double_negative(RS_106_io_sel_double_negative),
    .io_sel_double_positive(RS_106_io_sel_double_positive),
    .io_x(RS_106_io_x),
    .io_x_sub(RS_106_io_x_sub),
    .io_p(RS_106_io_p)
  );
  RS RS_107 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_107_io_sel_negative),
    .io_sel_positive(RS_107_io_sel_positive),
    .io_sel_double_negative(RS_107_io_sel_double_negative),
    .io_sel_double_positive(RS_107_io_sel_double_positive),
    .io_x(RS_107_io_x),
    .io_x_sub(RS_107_io_x_sub),
    .io_p(RS_107_io_p)
  );
  RS RS_108 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_108_io_sel_negative),
    .io_sel_positive(RS_108_io_sel_positive),
    .io_sel_double_negative(RS_108_io_sel_double_negative),
    .io_sel_double_positive(RS_108_io_sel_double_positive),
    .io_x(RS_108_io_x),
    .io_x_sub(RS_108_io_x_sub),
    .io_p(RS_108_io_p)
  );
  RS RS_109 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_109_io_sel_negative),
    .io_sel_positive(RS_109_io_sel_positive),
    .io_sel_double_negative(RS_109_io_sel_double_negative),
    .io_sel_double_positive(RS_109_io_sel_double_positive),
    .io_x(RS_109_io_x),
    .io_x_sub(RS_109_io_x_sub),
    .io_p(RS_109_io_p)
  );
  RS RS_110 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_110_io_sel_negative),
    .io_sel_positive(RS_110_io_sel_positive),
    .io_sel_double_negative(RS_110_io_sel_double_negative),
    .io_sel_double_positive(RS_110_io_sel_double_positive),
    .io_x(RS_110_io_x),
    .io_x_sub(RS_110_io_x_sub),
    .io_p(RS_110_io_p)
  );
  RS RS_111 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_111_io_sel_negative),
    .io_sel_positive(RS_111_io_sel_positive),
    .io_sel_double_negative(RS_111_io_sel_double_negative),
    .io_sel_double_positive(RS_111_io_sel_double_positive),
    .io_x(RS_111_io_x),
    .io_x_sub(RS_111_io_x_sub),
    .io_p(RS_111_io_p)
  );
  RS RS_112 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_112_io_sel_negative),
    .io_sel_positive(RS_112_io_sel_positive),
    .io_sel_double_negative(RS_112_io_sel_double_negative),
    .io_sel_double_positive(RS_112_io_sel_double_positive),
    .io_x(RS_112_io_x),
    .io_x_sub(RS_112_io_x_sub),
    .io_p(RS_112_io_p)
  );
  RS RS_113 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_113_io_sel_negative),
    .io_sel_positive(RS_113_io_sel_positive),
    .io_sel_double_negative(RS_113_io_sel_double_negative),
    .io_sel_double_positive(RS_113_io_sel_double_positive),
    .io_x(RS_113_io_x),
    .io_x_sub(RS_113_io_x_sub),
    .io_p(RS_113_io_p)
  );
  RS RS_114 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_114_io_sel_negative),
    .io_sel_positive(RS_114_io_sel_positive),
    .io_sel_double_negative(RS_114_io_sel_double_negative),
    .io_sel_double_positive(RS_114_io_sel_double_positive),
    .io_x(RS_114_io_x),
    .io_x_sub(RS_114_io_x_sub),
    .io_p(RS_114_io_p)
  );
  RS RS_115 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_115_io_sel_negative),
    .io_sel_positive(RS_115_io_sel_positive),
    .io_sel_double_negative(RS_115_io_sel_double_negative),
    .io_sel_double_positive(RS_115_io_sel_double_positive),
    .io_x(RS_115_io_x),
    .io_x_sub(RS_115_io_x_sub),
    .io_p(RS_115_io_p)
  );
  RS RS_116 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_116_io_sel_negative),
    .io_sel_positive(RS_116_io_sel_positive),
    .io_sel_double_negative(RS_116_io_sel_double_negative),
    .io_sel_double_positive(RS_116_io_sel_double_positive),
    .io_x(RS_116_io_x),
    .io_x_sub(RS_116_io_x_sub),
    .io_p(RS_116_io_p)
  );
  RS RS_117 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_117_io_sel_negative),
    .io_sel_positive(RS_117_io_sel_positive),
    .io_sel_double_negative(RS_117_io_sel_double_negative),
    .io_sel_double_positive(RS_117_io_sel_double_positive),
    .io_x(RS_117_io_x),
    .io_x_sub(RS_117_io_x_sub),
    .io_p(RS_117_io_p)
  );
  RS RS_118 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_118_io_sel_negative),
    .io_sel_positive(RS_118_io_sel_positive),
    .io_sel_double_negative(RS_118_io_sel_double_negative),
    .io_sel_double_positive(RS_118_io_sel_double_positive),
    .io_x(RS_118_io_x),
    .io_x_sub(RS_118_io_x_sub),
    .io_p(RS_118_io_p)
  );
  RS RS_119 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_119_io_sel_negative),
    .io_sel_positive(RS_119_io_sel_positive),
    .io_sel_double_negative(RS_119_io_sel_double_negative),
    .io_sel_double_positive(RS_119_io_sel_double_positive),
    .io_x(RS_119_io_x),
    .io_x_sub(RS_119_io_x_sub),
    .io_p(RS_119_io_p)
  );
  RS RS_120 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_120_io_sel_negative),
    .io_sel_positive(RS_120_io_sel_positive),
    .io_sel_double_negative(RS_120_io_sel_double_negative),
    .io_sel_double_positive(RS_120_io_sel_double_positive),
    .io_x(RS_120_io_x),
    .io_x_sub(RS_120_io_x_sub),
    .io_p(RS_120_io_p)
  );
  RS RS_121 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_121_io_sel_negative),
    .io_sel_positive(RS_121_io_sel_positive),
    .io_sel_double_negative(RS_121_io_sel_double_negative),
    .io_sel_double_positive(RS_121_io_sel_double_positive),
    .io_x(RS_121_io_x),
    .io_x_sub(RS_121_io_x_sub),
    .io_p(RS_121_io_p)
  );
  RS RS_122 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_122_io_sel_negative),
    .io_sel_positive(RS_122_io_sel_positive),
    .io_sel_double_negative(RS_122_io_sel_double_negative),
    .io_sel_double_positive(RS_122_io_sel_double_positive),
    .io_x(RS_122_io_x),
    .io_x_sub(RS_122_io_x_sub),
    .io_p(RS_122_io_p)
  );
  RS RS_123 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_123_io_sel_negative),
    .io_sel_positive(RS_123_io_sel_positive),
    .io_sel_double_negative(RS_123_io_sel_double_negative),
    .io_sel_double_positive(RS_123_io_sel_double_positive),
    .io_x(RS_123_io_x),
    .io_x_sub(RS_123_io_x_sub),
    .io_p(RS_123_io_p)
  );
  RS RS_124 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_124_io_sel_negative),
    .io_sel_positive(RS_124_io_sel_positive),
    .io_sel_double_negative(RS_124_io_sel_double_negative),
    .io_sel_double_positive(RS_124_io_sel_double_positive),
    .io_x(RS_124_io_x),
    .io_x_sub(RS_124_io_x_sub),
    .io_p(RS_124_io_p)
  );
  RS RS_125 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_125_io_sel_negative),
    .io_sel_positive(RS_125_io_sel_positive),
    .io_sel_double_negative(RS_125_io_sel_double_negative),
    .io_sel_double_positive(RS_125_io_sel_double_positive),
    .io_x(RS_125_io_x),
    .io_x_sub(RS_125_io_x_sub),
    .io_p(RS_125_io_p)
  );
  RS RS_126 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_126_io_sel_negative),
    .io_sel_positive(RS_126_io_sel_positive),
    .io_sel_double_negative(RS_126_io_sel_double_negative),
    .io_sel_double_positive(RS_126_io_sel_double_positive),
    .io_x(RS_126_io_x),
    .io_x_sub(RS_126_io_x_sub),
    .io_p(RS_126_io_p)
  );
  RS RS_127 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_127_io_sel_negative),
    .io_sel_positive(RS_127_io_sel_positive),
    .io_sel_double_negative(RS_127_io_sel_double_negative),
    .io_sel_double_positive(RS_127_io_sel_double_positive),
    .io_x(RS_127_io_x),
    .io_x_sub(RS_127_io_x_sub),
    .io_p(RS_127_io_p)
  );
  RS RS_128 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_128_io_sel_negative),
    .io_sel_positive(RS_128_io_sel_positive),
    .io_sel_double_negative(RS_128_io_sel_double_negative),
    .io_sel_double_positive(RS_128_io_sel_double_positive),
    .io_x(RS_128_io_x),
    .io_x_sub(RS_128_io_x_sub),
    .io_p(RS_128_io_p)
  );
  RS RS_129 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_129_io_sel_negative),
    .io_sel_positive(RS_129_io_sel_positive),
    .io_sel_double_negative(RS_129_io_sel_double_negative),
    .io_sel_double_positive(RS_129_io_sel_double_positive),
    .io_x(RS_129_io_x),
    .io_x_sub(RS_129_io_x_sub),
    .io_p(RS_129_io_p)
  );
  RS RS_130 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_130_io_sel_negative),
    .io_sel_positive(RS_130_io_sel_positive),
    .io_sel_double_negative(RS_130_io_sel_double_negative),
    .io_sel_double_positive(RS_130_io_sel_double_positive),
    .io_x(RS_130_io_x),
    .io_x_sub(RS_130_io_x_sub),
    .io_p(RS_130_io_p)
  );
  RS RS_131 ( // @[BOOTH_gen.scala 15:42]
    .io_sel_negative(RS_131_io_sel_negative),
    .io_sel_positive(RS_131_io_sel_positive),
    .io_sel_double_negative(RS_131_io_sel_double_negative),
    .io_sel_double_positive(RS_131_io_sel_double_positive),
    .io_x(RS_131_io_x),
    .io_x_sub(RS_131_io_x_sub),
    .io_p(RS_131_io_p)
  );
  BOOTH_S BOOTH_S ( // @[BOOTH_gen.scala 16:21]
    .io_sel_negative(BOOTH_S_io_sel_negative),
    .io_sel_positive(BOOTH_S_io_sel_positive),
    .io_sel_double_negative(BOOTH_S_io_sel_double_negative),
    .io_sel_double_positive(BOOTH_S_io_sel_double_positive),
    .io_src(BOOTH_S_io_src)
  );
  assign io_out = {io_out_hi,io_out_lo}; // @[Cat.scala 31:58]
  assign RS_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 22:23]
  assign RS_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 23:23]
  assign RS_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 24:30]
  assign RS_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 25:30]
  assign RS_io_x = io_x[0]; // @[BOOTH_gen.scala 20:16]
  assign RS_io_x_sub = 1'h0; // @[BOOTH_gen.scala 15:20 21:16]
  assign RS_1_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_1_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_1_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_1_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_1_io_x = io_x[1]; // @[BOOTH_gen.scala 28:20]
  assign RS_1_io_x_sub = io_x[0]; // @[BOOTH_gen.scala 29:24]
  assign RS_2_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_2_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_2_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_2_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_2_io_x = io_x[2]; // @[BOOTH_gen.scala 28:20]
  assign RS_2_io_x_sub = io_x[1]; // @[BOOTH_gen.scala 29:24]
  assign RS_3_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_3_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_3_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_3_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_3_io_x = io_x[3]; // @[BOOTH_gen.scala 28:20]
  assign RS_3_io_x_sub = io_x[2]; // @[BOOTH_gen.scala 29:24]
  assign RS_4_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_4_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_4_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_4_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_4_io_x = io_x[4]; // @[BOOTH_gen.scala 28:20]
  assign RS_4_io_x_sub = io_x[3]; // @[BOOTH_gen.scala 29:24]
  assign RS_5_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_5_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_5_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_5_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_5_io_x = io_x[5]; // @[BOOTH_gen.scala 28:20]
  assign RS_5_io_x_sub = io_x[4]; // @[BOOTH_gen.scala 29:24]
  assign RS_6_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_6_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_6_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_6_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_6_io_x = io_x[6]; // @[BOOTH_gen.scala 28:20]
  assign RS_6_io_x_sub = io_x[5]; // @[BOOTH_gen.scala 29:24]
  assign RS_7_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_7_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_7_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_7_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_7_io_x = io_x[7]; // @[BOOTH_gen.scala 28:20]
  assign RS_7_io_x_sub = io_x[6]; // @[BOOTH_gen.scala 29:24]
  assign RS_8_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_8_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_8_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_8_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_8_io_x = io_x[8]; // @[BOOTH_gen.scala 28:20]
  assign RS_8_io_x_sub = io_x[7]; // @[BOOTH_gen.scala 29:24]
  assign RS_9_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_9_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_9_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_9_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_9_io_x = io_x[9]; // @[BOOTH_gen.scala 28:20]
  assign RS_9_io_x_sub = io_x[8]; // @[BOOTH_gen.scala 29:24]
  assign RS_10_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_10_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_10_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_10_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_10_io_x = io_x[10]; // @[BOOTH_gen.scala 28:20]
  assign RS_10_io_x_sub = io_x[9]; // @[BOOTH_gen.scala 29:24]
  assign RS_11_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_11_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_11_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_11_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_11_io_x = io_x[11]; // @[BOOTH_gen.scala 28:20]
  assign RS_11_io_x_sub = io_x[10]; // @[BOOTH_gen.scala 29:24]
  assign RS_12_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_12_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_12_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_12_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_12_io_x = io_x[12]; // @[BOOTH_gen.scala 28:20]
  assign RS_12_io_x_sub = io_x[11]; // @[BOOTH_gen.scala 29:24]
  assign RS_13_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_13_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_13_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_13_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_13_io_x = io_x[13]; // @[BOOTH_gen.scala 28:20]
  assign RS_13_io_x_sub = io_x[12]; // @[BOOTH_gen.scala 29:24]
  assign RS_14_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_14_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_14_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_14_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_14_io_x = io_x[14]; // @[BOOTH_gen.scala 28:20]
  assign RS_14_io_x_sub = io_x[13]; // @[BOOTH_gen.scala 29:24]
  assign RS_15_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_15_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_15_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_15_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_15_io_x = io_x[15]; // @[BOOTH_gen.scala 28:20]
  assign RS_15_io_x_sub = io_x[14]; // @[BOOTH_gen.scala 29:24]
  assign RS_16_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_16_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_16_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_16_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_16_io_x = io_x[16]; // @[BOOTH_gen.scala 28:20]
  assign RS_16_io_x_sub = io_x[15]; // @[BOOTH_gen.scala 29:24]
  assign RS_17_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_17_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_17_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_17_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_17_io_x = io_x[17]; // @[BOOTH_gen.scala 28:20]
  assign RS_17_io_x_sub = io_x[16]; // @[BOOTH_gen.scala 29:24]
  assign RS_18_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_18_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_18_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_18_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_18_io_x = io_x[18]; // @[BOOTH_gen.scala 28:20]
  assign RS_18_io_x_sub = io_x[17]; // @[BOOTH_gen.scala 29:24]
  assign RS_19_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_19_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_19_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_19_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_19_io_x = io_x[19]; // @[BOOTH_gen.scala 28:20]
  assign RS_19_io_x_sub = io_x[18]; // @[BOOTH_gen.scala 29:24]
  assign RS_20_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_20_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_20_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_20_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_20_io_x = io_x[20]; // @[BOOTH_gen.scala 28:20]
  assign RS_20_io_x_sub = io_x[19]; // @[BOOTH_gen.scala 29:24]
  assign RS_21_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_21_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_21_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_21_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_21_io_x = io_x[21]; // @[BOOTH_gen.scala 28:20]
  assign RS_21_io_x_sub = io_x[20]; // @[BOOTH_gen.scala 29:24]
  assign RS_22_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_22_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_22_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_22_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_22_io_x = io_x[22]; // @[BOOTH_gen.scala 28:20]
  assign RS_22_io_x_sub = io_x[21]; // @[BOOTH_gen.scala 29:24]
  assign RS_23_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_23_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_23_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_23_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_23_io_x = io_x[23]; // @[BOOTH_gen.scala 28:20]
  assign RS_23_io_x_sub = io_x[22]; // @[BOOTH_gen.scala 29:24]
  assign RS_24_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_24_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_24_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_24_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_24_io_x = io_x[24]; // @[BOOTH_gen.scala 28:20]
  assign RS_24_io_x_sub = io_x[23]; // @[BOOTH_gen.scala 29:24]
  assign RS_25_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_25_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_25_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_25_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_25_io_x = io_x[25]; // @[BOOTH_gen.scala 28:20]
  assign RS_25_io_x_sub = io_x[24]; // @[BOOTH_gen.scala 29:24]
  assign RS_26_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_26_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_26_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_26_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_26_io_x = io_x[26]; // @[BOOTH_gen.scala 28:20]
  assign RS_26_io_x_sub = io_x[25]; // @[BOOTH_gen.scala 29:24]
  assign RS_27_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_27_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_27_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_27_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_27_io_x = io_x[27]; // @[BOOTH_gen.scala 28:20]
  assign RS_27_io_x_sub = io_x[26]; // @[BOOTH_gen.scala 29:24]
  assign RS_28_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_28_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_28_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_28_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_28_io_x = io_x[28]; // @[BOOTH_gen.scala 28:20]
  assign RS_28_io_x_sub = io_x[27]; // @[BOOTH_gen.scala 29:24]
  assign RS_29_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_29_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_29_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_29_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_29_io_x = io_x[29]; // @[BOOTH_gen.scala 28:20]
  assign RS_29_io_x_sub = io_x[28]; // @[BOOTH_gen.scala 29:24]
  assign RS_30_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_30_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_30_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_30_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_30_io_x = io_x[30]; // @[BOOTH_gen.scala 28:20]
  assign RS_30_io_x_sub = io_x[29]; // @[BOOTH_gen.scala 29:24]
  assign RS_31_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_31_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_31_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_31_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_31_io_x = io_x[31]; // @[BOOTH_gen.scala 28:20]
  assign RS_31_io_x_sub = io_x[30]; // @[BOOTH_gen.scala 29:24]
  assign RS_32_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_32_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_32_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_32_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_32_io_x = io_x[32]; // @[BOOTH_gen.scala 28:20]
  assign RS_32_io_x_sub = io_x[31]; // @[BOOTH_gen.scala 29:24]
  assign RS_33_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_33_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_33_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_33_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_33_io_x = io_x[33]; // @[BOOTH_gen.scala 28:20]
  assign RS_33_io_x_sub = io_x[32]; // @[BOOTH_gen.scala 29:24]
  assign RS_34_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_34_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_34_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_34_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_34_io_x = io_x[34]; // @[BOOTH_gen.scala 28:20]
  assign RS_34_io_x_sub = io_x[33]; // @[BOOTH_gen.scala 29:24]
  assign RS_35_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_35_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_35_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_35_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_35_io_x = io_x[35]; // @[BOOTH_gen.scala 28:20]
  assign RS_35_io_x_sub = io_x[34]; // @[BOOTH_gen.scala 29:24]
  assign RS_36_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_36_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_36_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_36_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_36_io_x = io_x[36]; // @[BOOTH_gen.scala 28:20]
  assign RS_36_io_x_sub = io_x[35]; // @[BOOTH_gen.scala 29:24]
  assign RS_37_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_37_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_37_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_37_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_37_io_x = io_x[37]; // @[BOOTH_gen.scala 28:20]
  assign RS_37_io_x_sub = io_x[36]; // @[BOOTH_gen.scala 29:24]
  assign RS_38_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_38_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_38_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_38_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_38_io_x = io_x[38]; // @[BOOTH_gen.scala 28:20]
  assign RS_38_io_x_sub = io_x[37]; // @[BOOTH_gen.scala 29:24]
  assign RS_39_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_39_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_39_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_39_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_39_io_x = io_x[39]; // @[BOOTH_gen.scala 28:20]
  assign RS_39_io_x_sub = io_x[38]; // @[BOOTH_gen.scala 29:24]
  assign RS_40_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_40_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_40_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_40_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_40_io_x = io_x[40]; // @[BOOTH_gen.scala 28:20]
  assign RS_40_io_x_sub = io_x[39]; // @[BOOTH_gen.scala 29:24]
  assign RS_41_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_41_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_41_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_41_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_41_io_x = io_x[41]; // @[BOOTH_gen.scala 28:20]
  assign RS_41_io_x_sub = io_x[40]; // @[BOOTH_gen.scala 29:24]
  assign RS_42_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_42_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_42_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_42_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_42_io_x = io_x[42]; // @[BOOTH_gen.scala 28:20]
  assign RS_42_io_x_sub = io_x[41]; // @[BOOTH_gen.scala 29:24]
  assign RS_43_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_43_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_43_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_43_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_43_io_x = io_x[43]; // @[BOOTH_gen.scala 28:20]
  assign RS_43_io_x_sub = io_x[42]; // @[BOOTH_gen.scala 29:24]
  assign RS_44_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_44_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_44_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_44_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_44_io_x = io_x[44]; // @[BOOTH_gen.scala 28:20]
  assign RS_44_io_x_sub = io_x[43]; // @[BOOTH_gen.scala 29:24]
  assign RS_45_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_45_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_45_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_45_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_45_io_x = io_x[45]; // @[BOOTH_gen.scala 28:20]
  assign RS_45_io_x_sub = io_x[44]; // @[BOOTH_gen.scala 29:24]
  assign RS_46_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_46_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_46_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_46_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_46_io_x = io_x[46]; // @[BOOTH_gen.scala 28:20]
  assign RS_46_io_x_sub = io_x[45]; // @[BOOTH_gen.scala 29:24]
  assign RS_47_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_47_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_47_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_47_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_47_io_x = io_x[47]; // @[BOOTH_gen.scala 28:20]
  assign RS_47_io_x_sub = io_x[46]; // @[BOOTH_gen.scala 29:24]
  assign RS_48_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_48_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_48_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_48_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_48_io_x = io_x[48]; // @[BOOTH_gen.scala 28:20]
  assign RS_48_io_x_sub = io_x[47]; // @[BOOTH_gen.scala 29:24]
  assign RS_49_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_49_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_49_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_49_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_49_io_x = io_x[49]; // @[BOOTH_gen.scala 28:20]
  assign RS_49_io_x_sub = io_x[48]; // @[BOOTH_gen.scala 29:24]
  assign RS_50_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_50_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_50_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_50_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_50_io_x = io_x[50]; // @[BOOTH_gen.scala 28:20]
  assign RS_50_io_x_sub = io_x[49]; // @[BOOTH_gen.scala 29:24]
  assign RS_51_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_51_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_51_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_51_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_51_io_x = io_x[51]; // @[BOOTH_gen.scala 28:20]
  assign RS_51_io_x_sub = io_x[50]; // @[BOOTH_gen.scala 29:24]
  assign RS_52_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_52_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_52_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_52_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_52_io_x = io_x[52]; // @[BOOTH_gen.scala 28:20]
  assign RS_52_io_x_sub = io_x[51]; // @[BOOTH_gen.scala 29:24]
  assign RS_53_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_53_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_53_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_53_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_53_io_x = io_x[53]; // @[BOOTH_gen.scala 28:20]
  assign RS_53_io_x_sub = io_x[52]; // @[BOOTH_gen.scala 29:24]
  assign RS_54_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_54_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_54_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_54_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_54_io_x = io_x[54]; // @[BOOTH_gen.scala 28:20]
  assign RS_54_io_x_sub = io_x[53]; // @[BOOTH_gen.scala 29:24]
  assign RS_55_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_55_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_55_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_55_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_55_io_x = io_x[55]; // @[BOOTH_gen.scala 28:20]
  assign RS_55_io_x_sub = io_x[54]; // @[BOOTH_gen.scala 29:24]
  assign RS_56_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_56_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_56_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_56_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_56_io_x = io_x[56]; // @[BOOTH_gen.scala 28:20]
  assign RS_56_io_x_sub = io_x[55]; // @[BOOTH_gen.scala 29:24]
  assign RS_57_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_57_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_57_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_57_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_57_io_x = io_x[57]; // @[BOOTH_gen.scala 28:20]
  assign RS_57_io_x_sub = io_x[56]; // @[BOOTH_gen.scala 29:24]
  assign RS_58_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_58_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_58_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_58_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_58_io_x = io_x[58]; // @[BOOTH_gen.scala 28:20]
  assign RS_58_io_x_sub = io_x[57]; // @[BOOTH_gen.scala 29:24]
  assign RS_59_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_59_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_59_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_59_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_59_io_x = io_x[59]; // @[BOOTH_gen.scala 28:20]
  assign RS_59_io_x_sub = io_x[58]; // @[BOOTH_gen.scala 29:24]
  assign RS_60_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_60_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_60_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_60_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_60_io_x = io_x[60]; // @[BOOTH_gen.scala 28:20]
  assign RS_60_io_x_sub = io_x[59]; // @[BOOTH_gen.scala 29:24]
  assign RS_61_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_61_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_61_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_61_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_61_io_x = io_x[61]; // @[BOOTH_gen.scala 28:20]
  assign RS_61_io_x_sub = io_x[60]; // @[BOOTH_gen.scala 29:24]
  assign RS_62_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_62_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_62_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_62_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_62_io_x = io_x[62]; // @[BOOTH_gen.scala 28:20]
  assign RS_62_io_x_sub = io_x[61]; // @[BOOTH_gen.scala 29:24]
  assign RS_63_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_63_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_63_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_63_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_63_io_x = io_x[63]; // @[BOOTH_gen.scala 28:20]
  assign RS_63_io_x_sub = io_x[62]; // @[BOOTH_gen.scala 29:24]
  assign RS_64_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_64_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_64_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_64_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_64_io_x = io_x[64]; // @[BOOTH_gen.scala 28:20]
  assign RS_64_io_x_sub = io_x[63]; // @[BOOTH_gen.scala 29:24]
  assign RS_65_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_65_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_65_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_65_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_65_io_x = io_x[65]; // @[BOOTH_gen.scala 28:20]
  assign RS_65_io_x_sub = io_x[64]; // @[BOOTH_gen.scala 29:24]
  assign RS_66_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_66_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_66_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_66_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_66_io_x = io_x[66]; // @[BOOTH_gen.scala 28:20]
  assign RS_66_io_x_sub = io_x[65]; // @[BOOTH_gen.scala 29:24]
  assign RS_67_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_67_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_67_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_67_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_67_io_x = io_x[67]; // @[BOOTH_gen.scala 28:20]
  assign RS_67_io_x_sub = io_x[66]; // @[BOOTH_gen.scala 29:24]
  assign RS_68_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_68_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_68_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_68_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_68_io_x = io_x[68]; // @[BOOTH_gen.scala 28:20]
  assign RS_68_io_x_sub = io_x[67]; // @[BOOTH_gen.scala 29:24]
  assign RS_69_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_69_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_69_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_69_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_69_io_x = io_x[69]; // @[BOOTH_gen.scala 28:20]
  assign RS_69_io_x_sub = io_x[68]; // @[BOOTH_gen.scala 29:24]
  assign RS_70_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_70_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_70_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_70_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_70_io_x = io_x[70]; // @[BOOTH_gen.scala 28:20]
  assign RS_70_io_x_sub = io_x[69]; // @[BOOTH_gen.scala 29:24]
  assign RS_71_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_71_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_71_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_71_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_71_io_x = io_x[71]; // @[BOOTH_gen.scala 28:20]
  assign RS_71_io_x_sub = io_x[70]; // @[BOOTH_gen.scala 29:24]
  assign RS_72_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_72_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_72_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_72_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_72_io_x = io_x[72]; // @[BOOTH_gen.scala 28:20]
  assign RS_72_io_x_sub = io_x[71]; // @[BOOTH_gen.scala 29:24]
  assign RS_73_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_73_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_73_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_73_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_73_io_x = io_x[73]; // @[BOOTH_gen.scala 28:20]
  assign RS_73_io_x_sub = io_x[72]; // @[BOOTH_gen.scala 29:24]
  assign RS_74_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_74_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_74_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_74_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_74_io_x = io_x[74]; // @[BOOTH_gen.scala 28:20]
  assign RS_74_io_x_sub = io_x[73]; // @[BOOTH_gen.scala 29:24]
  assign RS_75_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_75_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_75_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_75_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_75_io_x = io_x[75]; // @[BOOTH_gen.scala 28:20]
  assign RS_75_io_x_sub = io_x[74]; // @[BOOTH_gen.scala 29:24]
  assign RS_76_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_76_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_76_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_76_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_76_io_x = io_x[76]; // @[BOOTH_gen.scala 28:20]
  assign RS_76_io_x_sub = io_x[75]; // @[BOOTH_gen.scala 29:24]
  assign RS_77_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_77_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_77_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_77_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_77_io_x = io_x[77]; // @[BOOTH_gen.scala 28:20]
  assign RS_77_io_x_sub = io_x[76]; // @[BOOTH_gen.scala 29:24]
  assign RS_78_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_78_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_78_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_78_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_78_io_x = io_x[78]; // @[BOOTH_gen.scala 28:20]
  assign RS_78_io_x_sub = io_x[77]; // @[BOOTH_gen.scala 29:24]
  assign RS_79_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_79_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_79_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_79_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_79_io_x = io_x[79]; // @[BOOTH_gen.scala 28:20]
  assign RS_79_io_x_sub = io_x[78]; // @[BOOTH_gen.scala 29:24]
  assign RS_80_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_80_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_80_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_80_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_80_io_x = io_x[80]; // @[BOOTH_gen.scala 28:20]
  assign RS_80_io_x_sub = io_x[79]; // @[BOOTH_gen.scala 29:24]
  assign RS_81_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_81_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_81_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_81_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_81_io_x = io_x[81]; // @[BOOTH_gen.scala 28:20]
  assign RS_81_io_x_sub = io_x[80]; // @[BOOTH_gen.scala 29:24]
  assign RS_82_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_82_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_82_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_82_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_82_io_x = io_x[82]; // @[BOOTH_gen.scala 28:20]
  assign RS_82_io_x_sub = io_x[81]; // @[BOOTH_gen.scala 29:24]
  assign RS_83_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_83_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_83_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_83_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_83_io_x = io_x[83]; // @[BOOTH_gen.scala 28:20]
  assign RS_83_io_x_sub = io_x[82]; // @[BOOTH_gen.scala 29:24]
  assign RS_84_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_84_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_84_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_84_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_84_io_x = io_x[84]; // @[BOOTH_gen.scala 28:20]
  assign RS_84_io_x_sub = io_x[83]; // @[BOOTH_gen.scala 29:24]
  assign RS_85_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_85_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_85_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_85_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_85_io_x = io_x[85]; // @[BOOTH_gen.scala 28:20]
  assign RS_85_io_x_sub = io_x[84]; // @[BOOTH_gen.scala 29:24]
  assign RS_86_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_86_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_86_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_86_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_86_io_x = io_x[86]; // @[BOOTH_gen.scala 28:20]
  assign RS_86_io_x_sub = io_x[85]; // @[BOOTH_gen.scala 29:24]
  assign RS_87_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_87_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_87_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_87_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_87_io_x = io_x[87]; // @[BOOTH_gen.scala 28:20]
  assign RS_87_io_x_sub = io_x[86]; // @[BOOTH_gen.scala 29:24]
  assign RS_88_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_88_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_88_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_88_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_88_io_x = io_x[88]; // @[BOOTH_gen.scala 28:20]
  assign RS_88_io_x_sub = io_x[87]; // @[BOOTH_gen.scala 29:24]
  assign RS_89_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_89_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_89_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_89_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_89_io_x = io_x[89]; // @[BOOTH_gen.scala 28:20]
  assign RS_89_io_x_sub = io_x[88]; // @[BOOTH_gen.scala 29:24]
  assign RS_90_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_90_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_90_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_90_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_90_io_x = io_x[90]; // @[BOOTH_gen.scala 28:20]
  assign RS_90_io_x_sub = io_x[89]; // @[BOOTH_gen.scala 29:24]
  assign RS_91_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_91_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_91_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_91_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_91_io_x = io_x[91]; // @[BOOTH_gen.scala 28:20]
  assign RS_91_io_x_sub = io_x[90]; // @[BOOTH_gen.scala 29:24]
  assign RS_92_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_92_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_92_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_92_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_92_io_x = io_x[92]; // @[BOOTH_gen.scala 28:20]
  assign RS_92_io_x_sub = io_x[91]; // @[BOOTH_gen.scala 29:24]
  assign RS_93_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_93_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_93_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_93_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_93_io_x = io_x[93]; // @[BOOTH_gen.scala 28:20]
  assign RS_93_io_x_sub = io_x[92]; // @[BOOTH_gen.scala 29:24]
  assign RS_94_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_94_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_94_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_94_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_94_io_x = io_x[94]; // @[BOOTH_gen.scala 28:20]
  assign RS_94_io_x_sub = io_x[93]; // @[BOOTH_gen.scala 29:24]
  assign RS_95_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_95_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_95_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_95_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_95_io_x = io_x[95]; // @[BOOTH_gen.scala 28:20]
  assign RS_95_io_x_sub = io_x[94]; // @[BOOTH_gen.scala 29:24]
  assign RS_96_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_96_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_96_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_96_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_96_io_x = io_x[96]; // @[BOOTH_gen.scala 28:20]
  assign RS_96_io_x_sub = io_x[95]; // @[BOOTH_gen.scala 29:24]
  assign RS_97_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_97_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_97_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_97_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_97_io_x = io_x[97]; // @[BOOTH_gen.scala 28:20]
  assign RS_97_io_x_sub = io_x[96]; // @[BOOTH_gen.scala 29:24]
  assign RS_98_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_98_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_98_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_98_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_98_io_x = io_x[98]; // @[BOOTH_gen.scala 28:20]
  assign RS_98_io_x_sub = io_x[97]; // @[BOOTH_gen.scala 29:24]
  assign RS_99_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_99_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_99_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_99_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_99_io_x = io_x[99]; // @[BOOTH_gen.scala 28:20]
  assign RS_99_io_x_sub = io_x[98]; // @[BOOTH_gen.scala 29:24]
  assign RS_100_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_100_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_100_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_100_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_100_io_x = io_x[100]; // @[BOOTH_gen.scala 28:20]
  assign RS_100_io_x_sub = io_x[99]; // @[BOOTH_gen.scala 29:24]
  assign RS_101_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_101_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_101_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_101_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_101_io_x = io_x[101]; // @[BOOTH_gen.scala 28:20]
  assign RS_101_io_x_sub = io_x[100]; // @[BOOTH_gen.scala 29:24]
  assign RS_102_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_102_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_102_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_102_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_102_io_x = io_x[102]; // @[BOOTH_gen.scala 28:20]
  assign RS_102_io_x_sub = io_x[101]; // @[BOOTH_gen.scala 29:24]
  assign RS_103_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_103_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_103_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_103_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_103_io_x = io_x[103]; // @[BOOTH_gen.scala 28:20]
  assign RS_103_io_x_sub = io_x[102]; // @[BOOTH_gen.scala 29:24]
  assign RS_104_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_104_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_104_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_104_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_104_io_x = io_x[104]; // @[BOOTH_gen.scala 28:20]
  assign RS_104_io_x_sub = io_x[103]; // @[BOOTH_gen.scala 29:24]
  assign RS_105_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_105_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_105_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_105_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_105_io_x = io_x[105]; // @[BOOTH_gen.scala 28:20]
  assign RS_105_io_x_sub = io_x[104]; // @[BOOTH_gen.scala 29:24]
  assign RS_106_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_106_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_106_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_106_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_106_io_x = io_x[106]; // @[BOOTH_gen.scala 28:20]
  assign RS_106_io_x_sub = io_x[105]; // @[BOOTH_gen.scala 29:24]
  assign RS_107_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_107_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_107_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_107_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_107_io_x = io_x[107]; // @[BOOTH_gen.scala 28:20]
  assign RS_107_io_x_sub = io_x[106]; // @[BOOTH_gen.scala 29:24]
  assign RS_108_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_108_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_108_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_108_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_108_io_x = io_x[108]; // @[BOOTH_gen.scala 28:20]
  assign RS_108_io_x_sub = io_x[107]; // @[BOOTH_gen.scala 29:24]
  assign RS_109_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_109_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_109_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_109_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_109_io_x = io_x[109]; // @[BOOTH_gen.scala 28:20]
  assign RS_109_io_x_sub = io_x[108]; // @[BOOTH_gen.scala 29:24]
  assign RS_110_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_110_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_110_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_110_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_110_io_x = io_x[110]; // @[BOOTH_gen.scala 28:20]
  assign RS_110_io_x_sub = io_x[109]; // @[BOOTH_gen.scala 29:24]
  assign RS_111_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_111_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_111_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_111_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_111_io_x = io_x[111]; // @[BOOTH_gen.scala 28:20]
  assign RS_111_io_x_sub = io_x[110]; // @[BOOTH_gen.scala 29:24]
  assign RS_112_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_112_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_112_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_112_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_112_io_x = io_x[112]; // @[BOOTH_gen.scala 28:20]
  assign RS_112_io_x_sub = io_x[111]; // @[BOOTH_gen.scala 29:24]
  assign RS_113_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_113_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_113_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_113_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_113_io_x = io_x[113]; // @[BOOTH_gen.scala 28:20]
  assign RS_113_io_x_sub = io_x[112]; // @[BOOTH_gen.scala 29:24]
  assign RS_114_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_114_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_114_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_114_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_114_io_x = io_x[114]; // @[BOOTH_gen.scala 28:20]
  assign RS_114_io_x_sub = io_x[113]; // @[BOOTH_gen.scala 29:24]
  assign RS_115_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_115_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_115_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_115_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_115_io_x = io_x[115]; // @[BOOTH_gen.scala 28:20]
  assign RS_115_io_x_sub = io_x[114]; // @[BOOTH_gen.scala 29:24]
  assign RS_116_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_116_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_116_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_116_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_116_io_x = io_x[116]; // @[BOOTH_gen.scala 28:20]
  assign RS_116_io_x_sub = io_x[115]; // @[BOOTH_gen.scala 29:24]
  assign RS_117_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_117_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_117_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_117_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_117_io_x = io_x[117]; // @[BOOTH_gen.scala 28:20]
  assign RS_117_io_x_sub = io_x[116]; // @[BOOTH_gen.scala 29:24]
  assign RS_118_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_118_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_118_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_118_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_118_io_x = io_x[118]; // @[BOOTH_gen.scala 28:20]
  assign RS_118_io_x_sub = io_x[117]; // @[BOOTH_gen.scala 29:24]
  assign RS_119_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_119_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_119_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_119_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_119_io_x = io_x[119]; // @[BOOTH_gen.scala 28:20]
  assign RS_119_io_x_sub = io_x[118]; // @[BOOTH_gen.scala 29:24]
  assign RS_120_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_120_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_120_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_120_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_120_io_x = io_x[120]; // @[BOOTH_gen.scala 28:20]
  assign RS_120_io_x_sub = io_x[119]; // @[BOOTH_gen.scala 29:24]
  assign RS_121_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_121_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_121_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_121_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_121_io_x = io_x[121]; // @[BOOTH_gen.scala 28:20]
  assign RS_121_io_x_sub = io_x[120]; // @[BOOTH_gen.scala 29:24]
  assign RS_122_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_122_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_122_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_122_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_122_io_x = io_x[122]; // @[BOOTH_gen.scala 28:20]
  assign RS_122_io_x_sub = io_x[121]; // @[BOOTH_gen.scala 29:24]
  assign RS_123_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_123_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_123_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_123_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_123_io_x = io_x[123]; // @[BOOTH_gen.scala 28:20]
  assign RS_123_io_x_sub = io_x[122]; // @[BOOTH_gen.scala 29:24]
  assign RS_124_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_124_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_124_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_124_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_124_io_x = io_x[124]; // @[BOOTH_gen.scala 28:20]
  assign RS_124_io_x_sub = io_x[123]; // @[BOOTH_gen.scala 29:24]
  assign RS_125_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_125_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_125_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_125_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_125_io_x = io_x[125]; // @[BOOTH_gen.scala 28:20]
  assign RS_125_io_x_sub = io_x[124]; // @[BOOTH_gen.scala 29:24]
  assign RS_126_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_126_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_126_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_126_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_126_io_x = io_x[126]; // @[BOOTH_gen.scala 28:20]
  assign RS_126_io_x_sub = io_x[125]; // @[BOOTH_gen.scala 29:24]
  assign RS_127_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_127_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_127_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_127_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_127_io_x = io_x[127]; // @[BOOTH_gen.scala 28:20]
  assign RS_127_io_x_sub = io_x[126]; // @[BOOTH_gen.scala 29:24]
  assign RS_128_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_128_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_128_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_128_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_128_io_x = io_x[128]; // @[BOOTH_gen.scala 28:20]
  assign RS_128_io_x_sub = io_x[127]; // @[BOOTH_gen.scala 29:24]
  assign RS_129_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_129_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_129_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_129_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_129_io_x = io_x[129]; // @[BOOTH_gen.scala 28:20]
  assign RS_129_io_x_sub = io_x[128]; // @[BOOTH_gen.scala 29:24]
  assign RS_130_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_130_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_130_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_130_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_130_io_x = io_x[130]; // @[BOOTH_gen.scala 28:20]
  assign RS_130_io_x_sub = io_x[129]; // @[BOOTH_gen.scala 29:24]
  assign RS_131_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 15:20 30:27]
  assign RS_131_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 15:20 31:27]
  assign RS_131_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 15:20 32:34]
  assign RS_131_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 15:20 33:34]
  assign RS_131_io_x = io_x[131]; // @[BOOTH_gen.scala 28:20]
  assign RS_131_io_x_sub = io_x[130]; // @[BOOTH_gen.scala 29:24]
  assign BOOTH_S_io_src = io_y; // @[BOOTH_gen.scala 18:11]
endmodule
module MUL(
  input         clock,
  input         reset,
  input         io_mul_valid,
  input         io_flush,
  input         io_mulw,
  input  [1:0]  io_mul_signed,
  input  [63:0] io_multiplicand,
  input  [63:0] io_multiplier,
  output        io_mul_ready,
  output        io_out_valid,
  output [63:0] io_result_hi,
  output [63:0] io_result_lo
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire [131:0] BOOTH_gen_io_x; // @[MUL.scala 96:18]
  wire [2:0] BOOTH_gen_io_y; // @[MUL.scala 96:18]
  wire [131:0] BOOTH_gen_io_out; // @[MUL.scala 96:18]
  wire [65:0] multiplier = {io_mul_signed[1],io_multiplier,1'h0}; // @[Cat.scala 31:58]
  wire [65:0] multiplicand = {io_mul_signed[0],io_multiplicand,1'h0}; // @[Cat.scala 31:58]
  reg [131:0] multiplicand_reg; // @[MUL.scala 74:33]
  reg [65:0] multiplier_reg; // @[MUL.scala 75:31]
  reg [131:0] result; // @[MUL.scala 76:23]
  reg  start; // @[MUL.scala 77:22]
  reg [5:0] time_; // @[MUL.scala 78:21]
  wire  _GEN_1 = io_mul_valid | start; // @[MUL.scala 80:21 82:12 77:22]
  wire [5:0] _time_T_2 = time_ + 6'h1; // @[MUL.scala 92:38]
  wire  _multiplier_reg_T_1 = ~start & io_mul_valid; // @[MUL.scala 93:43]
  wire [133:0] _multiplicand_reg_T_2 = {multiplicand_reg, 2'h0}; // @[MUL.scala 94:93]
  wire [133:0] _multiplicand_reg_T_3 = _multiplier_reg_T_1 ? {{68'd0}, multiplicand} : _multiplicand_reg_T_2; // @[MUL.scala 94:26]
  wire [131:0] _result_T_2 = result + BOOTH_gen_io_out; // @[MUL.scala 100:42]
  wire [133:0] _GEN_6 = reset ? 134'h0 : _multiplicand_reg_T_3; // @[MUL.scala 74:{33,33} 94:20]
  BOOTH_gen BOOTH_gen ( // @[MUL.scala 96:18]
    .io_x(BOOTH_gen_io_x),
    .io_y(BOOTH_gen_io_y),
    .io_out(BOOTH_gen_io_out)
  );
  assign io_mul_ready = time_ == 6'h21; // @[MUL.scala 86:13]
  assign io_out_valid = time_ == 6'h21; // @[MUL.scala 86:13]
  assign io_result_hi = result[127:64]; // @[MUL.scala 102:25]
  assign io_result_lo = result[63:0]; // @[MUL.scala 103:25]
  assign BOOTH_gen_io_x = multiplicand_reg; // @[MUL.scala 98:8]
  assign BOOTH_gen_io_y = multiplier_reg[2:0]; // @[MUL.scala 97:25]
  always @(posedge clock) begin
    multiplicand_reg <= _GEN_6[131:0]; // @[MUL.scala 74:{33,33} 94:20]
    if (reset) begin // @[MUL.scala 75:31]
      multiplier_reg <= 66'h0; // @[MUL.scala 75:31]
    end else if (~start & io_mul_valid) begin // @[MUL.scala 93:24]
      multiplier_reg <= multiplier;
    end else begin
      multiplier_reg <= {{2'd0}, multiplier_reg[65:2]};
    end
    if (reset) begin // @[MUL.scala 76:23]
      result <= 132'h0; // @[MUL.scala 76:23]
    end else if (start) begin // @[MUL.scala 100:16]
      result <= _result_T_2;
    end
    if (reset) begin // @[MUL.scala 77:22]
      start <= 1'h0; // @[MUL.scala 77:22]
    end else if (time_ == 6'h21) begin // @[MUL.scala 86:22]
      start <= 1'h0; // @[MUL.scala 90:11]
    end else begin
      start <= _GEN_1;
    end
    if (reset) begin // @[MUL.scala 78:21]
      time_ <= 6'h0; // @[MUL.scala 78:21]
    end else if (start) begin // @[MUL.scala 92:14]
      time_ <= _time_T_2;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  multiplicand_reg = _RAND_0[131:0];
  _RAND_1 = {3{`RANDOM}};
  multiplier_reg = _RAND_1[65:0];
  _RAND_2 = {5{`RANDOM}};
  result = _RAND_2[131:0];
  _RAND_3 = {1{`RANDOM}};
  start = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  time_ = _RAND_4[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
