module IFU(
  input         clock,
  input         reset,
  input         io_reset,
  output [31:0] io_fd_bus_inst,
  output [31:0] io_fd_bus_pc,
  input         io_ds_allowin,
  output        io_fs_to_ds_valid,
  input         io_br_bus_br_taken,
  input  [31:0] io_br_bus_br_target,
  input         io_br_bus_rawblock,
  input  [63:0] io_br_bus_csr_rdata,
  input         io_br_bus_eval,
  input         io_br_bus_mret,
  output        io_inst_sram_req,
  output [63:0] io_inst_sram_addr,
  input  [63:0] io_inst_sram_rdata,
  input         io_inst_sram_addr_ok,
  input         io_inst_sram_data_ok
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg  fs_valid; // @[IFU.scala 23:35]
  reg  mid_handshake_inst; // @[IFU.scala 28:35]
  reg  inst_valid; // @[IFU.scala 29:35]
  reg [31:0] fs_inst; // @[IFU.scala 30:35]
  reg [63:0] fs_pc; // @[IFU.scala 31:35]
  reg [63:0] next_pc_R; // @[IFU.scala 32:35]
  reg  br_taken_R; // @[IFU.scala 33:35]
  reg  ex_taken_R; // @[IFU.scala 34:35]
  wire  prefs_ready_go = io_inst_sram_req & io_inst_sram_addr_ok; // @[IFU.scala 39:39]
  wire [63:0] _nextpc_T_1 = io_br_bus_csr_rdata + 64'h4; // @[IFU.scala 76:61]
  wire [63:0] _seq_pc_T_1 = fs_pc + 64'h4; // @[IFU.scala 75:26]
  wire [31:0] seq_pc = _seq_pc_T_1[31:0]; // @[IFU.scala 47:29 75:17]
  wire [31:0] _nextpc_T_2 = io_br_bus_br_taken ? io_br_bus_br_target : seq_pc; // @[IFU.scala 76:71]
  wire [63:0] _nextpc_T_3 = io_br_bus_mret ? _nextpc_T_1 : {{32'd0}, _nextpc_T_2}; // @[IFU.scala 76:44]
  wire [63:0] _nextpc_T_4 = io_br_bus_eval ? io_br_bus_csr_rdata : _nextpc_T_3; // @[IFU.scala 76:23]
  wire [31:0] nextpc = _nextpc_T_4[31:0]; // @[IFU.scala 48:29 76:17]
  wire  fs_ready_go = io_inst_sram_data_ok | inst_valid; // @[IFU.scala 80:45]
  wire  _fs_allow_in_T_1 = fs_ready_go & io_ds_allowin; // @[IFU.scala 81:49]
  wire  fs_allow_in = ~fs_valid | fs_ready_go & io_ds_allowin; // @[IFU.scala 81:34]
  wire  _T_6 = ~prefs_ready_go; // @[IFU.scala 64:14]
  wire  _GEN_1 = ~prefs_ready_go & io_br_bus_br_taken | br_taken_R; // @[IFU.scala 64:71 65:16 33:35]
  wire  _GEN_3 = _T_6 & (io_br_bus_mret | io_br_bus_eval) | ex_taken_R; // @[IFU.scala 71:77 72:16 34:35]
  wire [63:0] _final_next_pc_T_1 = br_taken_R | ex_taken_R ? next_pc_R : {{32'd0}, nextpc}; // @[IFU.scala 77:23]
  wire  _to_fs_valid_T = ~io_reset; // @[IFU.scala 79:24]
  wire  to_fs_valid = ~io_reset & prefs_ready_go; // @[IFU.scala 79:34]
  wire [31:0] final_next_pc = _final_next_pc_T_1[31:0]; // @[IFU.scala 35:32 77:17]
  wire  _GEN_7 = fs_allow_in ? 1'h0 : mid_handshake_inst; // @[IFU.scala 96:27 97:24 28:35]
  wire  _GEN_8 = io_inst_sram_addr_ok & io_inst_sram_req & ~fs_allow_in | _GEN_7; // @[IFU.scala 94:72 95:24]
  wire  _T_20 = ~io_ds_allowin; // @[IFU.scala 102:38]
  wire  _GEN_10 = io_inst_sram_data_ok & ~io_ds_allowin | inst_valid; // @[IFU.scala 102:54 103:16 29:35]
  assign io_fd_bus_inst = inst_valid ? fs_inst : io_inst_sram_rdata[31:0]; // @[IFU.scala 36:25]
  assign io_fd_bus_pc = fs_pc[31:0]; // @[IFU.scala 37:19]
  assign io_fs_to_ds_valid = fs_valid & fs_ready_go & ~io_br_bus_br_taken; // @[IFU.scala 82:48]
  assign io_inst_sram_req = _to_fs_valid_T & fs_allow_in & ~io_br_bus_rawblock & ~mid_handshake_inst; // @[IFU.scala 106:72]
  assign io_inst_sram_addr = {{32'd0}, final_next_pc}; // @[IFU.scala 108:21]
  always @(posedge clock) begin
    if (reset) begin // @[IFU.scala 23:35]
      fs_valid <= 1'h0; // @[IFU.scala 23:35]
    end else if (fs_allow_in) begin // @[IFU.scala 84:21]
      fs_valid <= to_fs_valid; // @[IFU.scala 85:14]
    end
    if (reset) begin // @[IFU.scala 28:35]
      mid_handshake_inst <= 1'h0; // @[IFU.scala 28:35]
    end else if (io_inst_sram_data_ok) begin // @[IFU.scala 92:30]
      mid_handshake_inst <= 1'h0; // @[IFU.scala 93:24]
    end else begin
      mid_handshake_inst <= _GEN_8;
    end
    if (reset) begin // @[IFU.scala 29:35]
      inst_valid <= 1'h0; // @[IFU.scala 29:35]
    end else if (_fs_allow_in_T_1) begin // @[IFU.scala 100:38]
      inst_valid <= 1'h0; // @[IFU.scala 101:16]
    end else begin
      inst_valid <= _GEN_10;
    end
    if (reset) begin // @[IFU.scala 30:35]
      fs_inst <= 32'h0; // @[IFU.scala 30:35]
    end else if (fs_ready_go & _T_20 & io_inst_sram_data_ok) begin // @[IFU.scala 110:63]
      fs_inst <= io_inst_sram_rdata[31:0]; // @[IFU.scala 111:13]
    end
    if (reset) begin // @[IFU.scala 31:35]
      fs_pc <= 64'h80000000; // @[IFU.scala 31:35]
    end else if (fs_allow_in & io_inst_sram_addr_ok) begin // @[IFU.scala 88:45]
      fs_pc <= {{32'd0}, final_next_pc}; // @[IFU.scala 89:11]
    end
    if (reset) begin // @[IFU.scala 32:35]
      next_pc_R <= 64'h80000000; // @[IFU.scala 32:35]
    end else if (io_br_bus_br_taken | io_br_bus_mret | io_br_bus_eval) begin // @[IFU.scala 57:34]
      next_pc_R <= {{32'd0}, nextpc}; // @[IFU.scala 58:15]
    end
    if (reset) begin // @[IFU.scala 33:35]
      br_taken_R <= 1'h0; // @[IFU.scala 33:35]
    end else if (br_taken_R & io_inst_sram_req & io_inst_sram_addr_ok & fs_allow_in) begin // @[IFU.scala 61:79]
      br_taken_R <= 1'h0; // @[IFU.scala 62:16]
    end else begin
      br_taken_R <= _GEN_1;
    end
    if (reset) begin // @[IFU.scala 34:35]
      ex_taken_R <= 1'h0; // @[IFU.scala 34:35]
    end else if (ex_taken_R & io_inst_sram_req & io_inst_sram_addr_ok & fs_allow_in) begin // @[IFU.scala 68:79]
      ex_taken_R <= 1'h0; // @[IFU.scala 69:16]
    end else begin
      ex_taken_R <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fs_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  mid_handshake_inst = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inst_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  fs_inst = _RAND_3[31:0];
  _RAND_4 = {2{`RANDOM}};
  fs_pc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  next_pc_R = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  br_taken_R = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  ex_taken_R = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Registers(
  input         clock,
  input         io_wen,
  input  [63:0] io_wdata,
  output [63:0] io_rdata1,
  output [63:0] io_rdata2,
  input  [4:0]  io_rs1,
  input  [4:0]  io_rs2,
  input  [4:0]  io_waddr,
  output [63:0] io_regs_0,
  output [63:0] io_regs_1,
  output [63:0] io_regs_2,
  output [63:0] io_regs_3,
  output [63:0] io_regs_4,
  output [63:0] io_regs_5,
  output [63:0] io_regs_6,
  output [63:0] io_regs_7,
  output [63:0] io_regs_8,
  output [63:0] io_regs_9,
  output [63:0] io_regs_10,
  output [63:0] io_regs_11,
  output [63:0] io_regs_12,
  output [63:0] io_regs_13,
  output [63:0] io_regs_14,
  output [63:0] io_regs_15,
  output [63:0] io_regs_16,
  output [63:0] io_regs_17,
  output [63:0] io_regs_18,
  output [63:0] io_regs_19,
  output [63:0] io_regs_20,
  output [63:0] io_regs_21,
  output [63:0] io_regs_22,
  output [63:0] io_regs_23,
  output [63:0] io_regs_24,
  output [63:0] io_regs_25,
  output [63:0] io_regs_26,
  output [63:0] io_regs_27,
  output [63:0] io_regs_28,
  output [63:0] io_regs_29,
  output [63:0] io_regs_30,
  output [63:0] io_regs_31
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [63:0] registers [0:31]; // @[Registers.scala 22:22]
  wire  registers_io_rdata1_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_rdata1_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_rdata1_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_rdata2_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_rdata2_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_rdata2_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_reg17_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_reg17_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_reg17_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_MPORT_1_en; // @[Registers.scala 22:22]
  wire [4:0] registers_MPORT_1_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_MPORT_1_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_0_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_0_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_0_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_1_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_1_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_1_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_2_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_2_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_2_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_3_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_3_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_3_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_4_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_4_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_4_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_5_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_5_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_5_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_6_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_6_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_6_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_7_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_7_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_7_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_8_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_8_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_8_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_9_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_9_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_9_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_10_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_10_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_10_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_11_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_11_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_11_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_12_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_12_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_12_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_13_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_13_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_13_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_14_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_14_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_14_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_15_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_15_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_15_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_16_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_16_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_16_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_17_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_17_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_17_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_18_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_18_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_18_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_19_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_19_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_19_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_20_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_20_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_20_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_21_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_21_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_21_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_22_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_22_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_22_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_23_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_23_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_23_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_24_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_24_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_24_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_25_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_25_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_25_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_26_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_26_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_26_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_27_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_27_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_27_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_28_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_28_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_28_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_29_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_29_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_29_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_30_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_30_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_30_MPORT_data; // @[Registers.scala 22:22]
  wire  registers_io_regs_31_MPORT_en; // @[Registers.scala 22:22]
  wire [4:0] registers_io_regs_31_MPORT_addr; // @[Registers.scala 22:22]
  wire [63:0] registers_io_regs_31_MPORT_data; // @[Registers.scala 22:22]
  wire [63:0] registers_MPORT_data; // @[Registers.scala 22:22]
  wire [4:0] registers_MPORT_addr; // @[Registers.scala 22:22]
  wire  registers_MPORT_mask; // @[Registers.scala 22:22]
  wire  registers_MPORT_en; // @[Registers.scala 22:22]
  wire  _T_1 = io_wen & io_waddr != 5'h0; // @[Registers.scala 27:37]
  assign registers_io_rdata1_MPORT_en = 1'h1;
  assign registers_io_rdata1_MPORT_addr = io_rs1;
  assign registers_io_rdata1_MPORT_data = registers[registers_io_rdata1_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_rdata2_MPORT_en = 1'h1;
  assign registers_io_rdata2_MPORT_addr = io_rs2;
  assign registers_io_rdata2_MPORT_data = registers[registers_io_rdata2_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_reg17_MPORT_en = 1'h1;
  assign registers_io_reg17_MPORT_addr = 5'h11;
  assign registers_io_reg17_MPORT_data = registers[registers_io_reg17_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_MPORT_1_en = 1'h1;
  assign registers_MPORT_1_addr = io_waddr;
  assign registers_MPORT_1_data = registers[registers_MPORT_1_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_0_MPORT_en = 1'h1;
  assign registers_io_regs_0_MPORT_addr = 5'h0;
  assign registers_io_regs_0_MPORT_data = registers[registers_io_regs_0_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_1_MPORT_en = 1'h1;
  assign registers_io_regs_1_MPORT_addr = 5'h1;
  assign registers_io_regs_1_MPORT_data = registers[registers_io_regs_1_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_2_MPORT_en = 1'h1;
  assign registers_io_regs_2_MPORT_addr = 5'h2;
  assign registers_io_regs_2_MPORT_data = registers[registers_io_regs_2_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_3_MPORT_en = 1'h1;
  assign registers_io_regs_3_MPORT_addr = 5'h3;
  assign registers_io_regs_3_MPORT_data = registers[registers_io_regs_3_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_4_MPORT_en = 1'h1;
  assign registers_io_regs_4_MPORT_addr = 5'h4;
  assign registers_io_regs_4_MPORT_data = registers[registers_io_regs_4_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_5_MPORT_en = 1'h1;
  assign registers_io_regs_5_MPORT_addr = 5'h5;
  assign registers_io_regs_5_MPORT_data = registers[registers_io_regs_5_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_6_MPORT_en = 1'h1;
  assign registers_io_regs_6_MPORT_addr = 5'h6;
  assign registers_io_regs_6_MPORT_data = registers[registers_io_regs_6_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_7_MPORT_en = 1'h1;
  assign registers_io_regs_7_MPORT_addr = 5'h7;
  assign registers_io_regs_7_MPORT_data = registers[registers_io_regs_7_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_8_MPORT_en = 1'h1;
  assign registers_io_regs_8_MPORT_addr = 5'h8;
  assign registers_io_regs_8_MPORT_data = registers[registers_io_regs_8_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_9_MPORT_en = 1'h1;
  assign registers_io_regs_9_MPORT_addr = 5'h9;
  assign registers_io_regs_9_MPORT_data = registers[registers_io_regs_9_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_10_MPORT_en = 1'h1;
  assign registers_io_regs_10_MPORT_addr = 5'ha;
  assign registers_io_regs_10_MPORT_data = registers[registers_io_regs_10_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_11_MPORT_en = 1'h1;
  assign registers_io_regs_11_MPORT_addr = 5'hb;
  assign registers_io_regs_11_MPORT_data = registers[registers_io_regs_11_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_12_MPORT_en = 1'h1;
  assign registers_io_regs_12_MPORT_addr = 5'hc;
  assign registers_io_regs_12_MPORT_data = registers[registers_io_regs_12_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_13_MPORT_en = 1'h1;
  assign registers_io_regs_13_MPORT_addr = 5'hd;
  assign registers_io_regs_13_MPORT_data = registers[registers_io_regs_13_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_14_MPORT_en = 1'h1;
  assign registers_io_regs_14_MPORT_addr = 5'he;
  assign registers_io_regs_14_MPORT_data = registers[registers_io_regs_14_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_15_MPORT_en = 1'h1;
  assign registers_io_regs_15_MPORT_addr = 5'hf;
  assign registers_io_regs_15_MPORT_data = registers[registers_io_regs_15_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_16_MPORT_en = 1'h1;
  assign registers_io_regs_16_MPORT_addr = 5'h10;
  assign registers_io_regs_16_MPORT_data = registers[registers_io_regs_16_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_17_MPORT_en = 1'h1;
  assign registers_io_regs_17_MPORT_addr = 5'h11;
  assign registers_io_regs_17_MPORT_data = registers[registers_io_regs_17_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_18_MPORT_en = 1'h1;
  assign registers_io_regs_18_MPORT_addr = 5'h12;
  assign registers_io_regs_18_MPORT_data = registers[registers_io_regs_18_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_19_MPORT_en = 1'h1;
  assign registers_io_regs_19_MPORT_addr = 5'h13;
  assign registers_io_regs_19_MPORT_data = registers[registers_io_regs_19_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_20_MPORT_en = 1'h1;
  assign registers_io_regs_20_MPORT_addr = 5'h14;
  assign registers_io_regs_20_MPORT_data = registers[registers_io_regs_20_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_21_MPORT_en = 1'h1;
  assign registers_io_regs_21_MPORT_addr = 5'h15;
  assign registers_io_regs_21_MPORT_data = registers[registers_io_regs_21_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_22_MPORT_en = 1'h1;
  assign registers_io_regs_22_MPORT_addr = 5'h16;
  assign registers_io_regs_22_MPORT_data = registers[registers_io_regs_22_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_23_MPORT_en = 1'h1;
  assign registers_io_regs_23_MPORT_addr = 5'h17;
  assign registers_io_regs_23_MPORT_data = registers[registers_io_regs_23_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_24_MPORT_en = 1'h1;
  assign registers_io_regs_24_MPORT_addr = 5'h18;
  assign registers_io_regs_24_MPORT_data = registers[registers_io_regs_24_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_25_MPORT_en = 1'h1;
  assign registers_io_regs_25_MPORT_addr = 5'h19;
  assign registers_io_regs_25_MPORT_data = registers[registers_io_regs_25_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_26_MPORT_en = 1'h1;
  assign registers_io_regs_26_MPORT_addr = 5'h1a;
  assign registers_io_regs_26_MPORT_data = registers[registers_io_regs_26_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_27_MPORT_en = 1'h1;
  assign registers_io_regs_27_MPORT_addr = 5'h1b;
  assign registers_io_regs_27_MPORT_data = registers[registers_io_regs_27_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_28_MPORT_en = 1'h1;
  assign registers_io_regs_28_MPORT_addr = 5'h1c;
  assign registers_io_regs_28_MPORT_data = registers[registers_io_regs_28_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_29_MPORT_en = 1'h1;
  assign registers_io_regs_29_MPORT_addr = 5'h1d;
  assign registers_io_regs_29_MPORT_data = registers[registers_io_regs_29_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_30_MPORT_en = 1'h1;
  assign registers_io_regs_30_MPORT_addr = 5'h1e;
  assign registers_io_regs_30_MPORT_data = registers[registers_io_regs_30_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_io_regs_31_MPORT_en = 1'h1;
  assign registers_io_regs_31_MPORT_addr = 5'h1f;
  assign registers_io_regs_31_MPORT_data = registers[registers_io_regs_31_MPORT_addr]; // @[Registers.scala 22:22]
  assign registers_MPORT_data = _T_1 ? io_wdata : registers_MPORT_1_data;
  assign registers_MPORT_addr = io_waddr;
  assign registers_MPORT_mask = 1'h1;
  assign registers_MPORT_en = 1'h1;
  assign io_rdata1 = io_rs1 == 5'h0 ? 64'h0 : registers_io_rdata1_MPORT_data; // @[Registers.scala 23:19]
  assign io_rdata2 = io_rs2 == 5'h0 ? 64'h0 : registers_io_rdata2_MPORT_data; // @[Registers.scala 24:19]
  assign io_regs_0 = registers_io_regs_0_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_1 = registers_io_regs_1_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_2 = registers_io_regs_2_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_3 = registers_io_regs_3_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_4 = registers_io_regs_4_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_5 = registers_io_regs_5_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_6 = registers_io_regs_6_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_7 = registers_io_regs_7_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_8 = registers_io_regs_8_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_9 = registers_io_regs_9_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_10 = registers_io_regs_10_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_11 = registers_io_regs_11_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_12 = registers_io_regs_12_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_13 = registers_io_regs_13_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_14 = registers_io_regs_14_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_15 = registers_io_regs_15_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_16 = registers_io_regs_16_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_17 = registers_io_regs_17_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_18 = registers_io_regs_18_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_19 = registers_io_regs_19_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_20 = registers_io_regs_20_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_21 = registers_io_regs_21_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_22 = registers_io_regs_22_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_23 = registers_io_regs_23_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_24 = registers_io_regs_24_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_25 = registers_io_regs_25_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_26 = registers_io_regs_26_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_27 = registers_io_regs_27_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_28 = registers_io_regs_28_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_29 = registers_io_regs_29_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_30 = registers_io_regs_30_MPORT_data; // @[Registers.scala 29:40]
  assign io_regs_31 = registers_io_regs_31_MPORT_data; // @[Registers.scala 29:40]
  always @(posedge clock) begin
    if (registers_MPORT_en & registers_MPORT_mask) begin
      registers[registers_MPORT_addr] <= registers_MPORT_data; // @[Registers.scala 22:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    registers[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CSR(
  input         clock,
  input         io_wen,
  input         io_ren,
  input  [63:0] io_wdata1,
  input  [63:0] io_wdata2,
  output [63:0] io_rdata,
  input  [4:0]  io_waddr1,
  input  [4:0]  io_waddr2,
  input  [4:0]  io_raddr,
  output [63:0] io_csrs_0,
  output [63:0] io_csrs_1,
  output [63:0] io_csrs_2,
  output [63:0] io_csrs_3,
  output [63:0] io_csrs_4
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
  reg [63:0] csr [0:4]; // @[CSR.scala 21:16]
  wire  csr_io_rdata_MPORT_en; // @[CSR.scala 21:16]
  wire [2:0] csr_io_rdata_MPORT_addr; // @[CSR.scala 21:16]
  wire [63:0] csr_io_rdata_MPORT_data; // @[CSR.scala 21:16]
  wire  csr_MPORT_1_en; // @[CSR.scala 21:16]
  wire [2:0] csr_MPORT_1_addr; // @[CSR.scala 21:16]
  wire [63:0] csr_MPORT_1_data; // @[CSR.scala 21:16]
  wire  csr_MPORT_3_en; // @[CSR.scala 21:16]
  wire [2:0] csr_MPORT_3_addr; // @[CSR.scala 21:16]
  wire [63:0] csr_MPORT_3_data; // @[CSR.scala 21:16]
  wire  csr_io_csrs_0_MPORT_en; // @[CSR.scala 21:16]
  wire [2:0] csr_io_csrs_0_MPORT_addr; // @[CSR.scala 21:16]
  wire [63:0] csr_io_csrs_0_MPORT_data; // @[CSR.scala 21:16]
  wire  csr_io_csrs_1_MPORT_en; // @[CSR.scala 21:16]
  wire [2:0] csr_io_csrs_1_MPORT_addr; // @[CSR.scala 21:16]
  wire [63:0] csr_io_csrs_1_MPORT_data; // @[CSR.scala 21:16]
  wire  csr_io_csrs_2_MPORT_en; // @[CSR.scala 21:16]
  wire [2:0] csr_io_csrs_2_MPORT_addr; // @[CSR.scala 21:16]
  wire [63:0] csr_io_csrs_2_MPORT_data; // @[CSR.scala 21:16]
  wire  csr_io_csrs_3_MPORT_en; // @[CSR.scala 21:16]
  wire [2:0] csr_io_csrs_3_MPORT_addr; // @[CSR.scala 21:16]
  wire [63:0] csr_io_csrs_3_MPORT_data; // @[CSR.scala 21:16]
  wire  csr_io_csrs_4_MPORT_en; // @[CSR.scala 21:16]
  wire [2:0] csr_io_csrs_4_MPORT_addr; // @[CSR.scala 21:16]
  wire [63:0] csr_io_csrs_4_MPORT_data; // @[CSR.scala 21:16]
  wire [63:0] csr_MPORT_data; // @[CSR.scala 21:16]
  wire [2:0] csr_MPORT_addr; // @[CSR.scala 21:16]
  wire  csr_MPORT_mask; // @[CSR.scala 21:16]
  wire  csr_MPORT_en; // @[CSR.scala 21:16]
  wire [63:0] csr_MPORT_2_data; // @[CSR.scala 21:16]
  wire [2:0] csr_MPORT_2_addr; // @[CSR.scala 21:16]
  wire  csr_MPORT_2_mask; // @[CSR.scala 21:16]
  wire  csr_MPORT_2_en; // @[CSR.scala 21:16]
  wire  _T_2 = io_wen & io_waddr1 != 5'h0; // @[CSR.scala 24:32]
  wire  _T_7 = io_wen & io_waddr2 != 5'h0; // @[CSR.scala 25:32]
  assign csr_io_rdata_MPORT_en = 1'h1;
  assign csr_io_rdata_MPORT_addr = io_raddr[2:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign csr_io_rdata_MPORT_data = csr[csr_io_rdata_MPORT_addr]; // @[CSR.scala 21:16]
  `else
  assign csr_io_rdata_MPORT_data = csr_io_rdata_MPORT_addr >= 3'h5 ? _RAND_1[63:0] : csr[csr_io_rdata_MPORT_addr]; // @[CSR.scala 21:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign csr_MPORT_1_en = 1'h1;
  assign csr_MPORT_1_addr = io_waddr1[2:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign csr_MPORT_1_data = csr[csr_MPORT_1_addr]; // @[CSR.scala 21:16]
  `else
  assign csr_MPORT_1_data = csr_MPORT_1_addr >= 3'h5 ? _RAND_2[63:0] : csr[csr_MPORT_1_addr]; // @[CSR.scala 21:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign csr_MPORT_3_en = 1'h1;
  assign csr_MPORT_3_addr = io_waddr2[2:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign csr_MPORT_3_data = csr[csr_MPORT_3_addr]; // @[CSR.scala 21:16]
  `else
  assign csr_MPORT_3_data = csr_MPORT_3_addr >= 3'h5 ? _RAND_3[63:0] : csr[csr_MPORT_3_addr]; // @[CSR.scala 21:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign csr_io_csrs_0_MPORT_en = 1'h1;
  assign csr_io_csrs_0_MPORT_addr = 3'h0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign csr_io_csrs_0_MPORT_data = csr[csr_io_csrs_0_MPORT_addr]; // @[CSR.scala 21:16]
  `else
  assign csr_io_csrs_0_MPORT_data = csr_io_csrs_0_MPORT_addr >= 3'h5 ? _RAND_4[63:0] : csr[csr_io_csrs_0_MPORT_addr]; // @[CSR.scala 21:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign csr_io_csrs_1_MPORT_en = 1'h1;
  assign csr_io_csrs_1_MPORT_addr = 3'h1;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign csr_io_csrs_1_MPORT_data = csr[csr_io_csrs_1_MPORT_addr]; // @[CSR.scala 21:16]
  `else
  assign csr_io_csrs_1_MPORT_data = csr_io_csrs_1_MPORT_addr >= 3'h5 ? _RAND_5[63:0] : csr[csr_io_csrs_1_MPORT_addr]; // @[CSR.scala 21:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign csr_io_csrs_2_MPORT_en = 1'h1;
  assign csr_io_csrs_2_MPORT_addr = 3'h2;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign csr_io_csrs_2_MPORT_data = csr[csr_io_csrs_2_MPORT_addr]; // @[CSR.scala 21:16]
  `else
  assign csr_io_csrs_2_MPORT_data = csr_io_csrs_2_MPORT_addr >= 3'h5 ? _RAND_6[63:0] : csr[csr_io_csrs_2_MPORT_addr]; // @[CSR.scala 21:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign csr_io_csrs_3_MPORT_en = 1'h1;
  assign csr_io_csrs_3_MPORT_addr = 3'h3;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign csr_io_csrs_3_MPORT_data = csr[csr_io_csrs_3_MPORT_addr]; // @[CSR.scala 21:16]
  `else
  assign csr_io_csrs_3_MPORT_data = csr_io_csrs_3_MPORT_addr >= 3'h5 ? _RAND_7[63:0] : csr[csr_io_csrs_3_MPORT_addr]; // @[CSR.scala 21:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign csr_io_csrs_4_MPORT_en = 1'h1;
  assign csr_io_csrs_4_MPORT_addr = 3'h4;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign csr_io_csrs_4_MPORT_data = csr[csr_io_csrs_4_MPORT_addr]; // @[CSR.scala 21:16]
  `else
  assign csr_io_csrs_4_MPORT_data = csr_io_csrs_4_MPORT_addr >= 3'h5 ? _RAND_8[63:0] : csr[csr_io_csrs_4_MPORT_addr]; // @[CSR.scala 21:16]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign csr_MPORT_data = _T_2 ? io_wdata1 : csr_MPORT_1_data;
  assign csr_MPORT_addr = io_waddr1[2:0];
  assign csr_MPORT_mask = 1'h1;
  assign csr_MPORT_en = 1'h1;
  assign csr_MPORT_2_data = _T_7 ? io_wdata2 : csr_MPORT_3_data;
  assign csr_MPORT_2_addr = io_waddr2[2:0];
  assign csr_MPORT_2_mask = 1'h1;
  assign csr_MPORT_2_en = 1'h1;
  assign io_rdata = io_ren ? csr_io_rdata_MPORT_data : 64'h0; // @[CSR.scala 22:18]
  assign io_csrs_0 = csr_io_csrs_0_MPORT_data; // @[CSR.scala 27:39]
  assign io_csrs_1 = csr_io_csrs_1_MPORT_data; // @[CSR.scala 27:39]
  assign io_csrs_2 = csr_io_csrs_2_MPORT_data; // @[CSR.scala 27:39]
  assign io_csrs_3 = csr_io_csrs_3_MPORT_data; // @[CSR.scala 27:39]
  assign io_csrs_4 = csr_io_csrs_4_MPORT_data; // @[CSR.scala 27:39]
  always @(posedge clock) begin
    if (csr_MPORT_en & csr_MPORT_mask) begin
      csr[csr_MPORT_addr] <= csr_MPORT_data; // @[CSR.scala 21:16]
    end
    if (csr_MPORT_2_en & csr_MPORT_2_mask) begin
      csr[csr_MPORT_2_addr] <= csr_MPORT_2_data; // @[CSR.scala 21:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {2{`RANDOM}};
  _RAND_2 = {2{`RANDOM}};
  _RAND_3 = {2{`RANDOM}};
  _RAND_4 = {2{`RANDOM}};
  _RAND_5 = {2{`RANDOM}};
  _RAND_6 = {2{`RANDOM}};
  _RAND_7 = {2{`RANDOM}};
  _RAND_8 = {2{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 5; initvar = initvar+1)
    csr[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IDU(
  input         clock,
  input         reset,
  input         io_es_allowin,
  output        io_ds_allowin,
  input         io_fs_to_ds_valid,
  output        io_ds_to_es_valid,
  input  [31:0] io_fd_bus_inst,
  input  [31:0] io_fd_bus_pc,
  output [7:0]  io_de_bus_OP,
  output        io_de_bus_res_from_mem,
  output        io_de_bus_gr_we,
  output        io_de_bus_MemWen,
  output [7:0]  io_de_bus_wmask,
  output [31:0] io_de_bus_ds_pc,
  output [4:0]  io_de_bus_dest,
  output [63:0] io_de_bus_imm,
  output [63:0] io_de_bus_rdata1,
  output [63:0] io_de_bus_rdata2,
  output [2:0]  io_de_bus_ld_type,
  output [31:0] io_de_bus_inst,
  output [63:0] io_de_bus_csr_rdata,
  output [2:0]  io_de_bus_csr_waddr1,
  output [2:0]  io_de_bus_csr_waddr2,
  output [2:0]  io_de_bus_csr_raddr,
  output        io_de_bus_csr_ren,
  output        io_de_bus_csr_wen,
  output        io_de_bus_eval,
  output        io_de_bus_is_ld,
  output        io_br_bus_br_taken,
  output [31:0] io_br_bus_br_target,
  output        io_br_bus_rawblock,
  output [63:0] io_br_bus_csr_rdata,
  output        io_br_bus_eval,
  output        io_br_bus_mret,
  input         io_rf_bus_rf_we,
  input  [4:0]  io_rf_bus_rf_waddr,
  input  [63:0] io_rf_bus_rf_wdata,
  input  [31:0] io_rf_bus_wb_pc,
  input  [31:0] io_rf_bus_wb_inst,
  input  [63:0] io_rf_bus_csr_wdata,
  input         io_rf_bus_csr_wen,
  input  [2:0]  io_rf_bus_csr_waddr1,
  input  [2:0]  io_rf_bus_csr_waddr2,
  input         io_rf_bus_eval,
  input         io_es_dest_valid_gr_we,
  input         io_es_dest_valid_es_valid,
  input  [4:0]  io_es_dest_valid_dest,
  input  [63:0] io_es_dest_valid_es_forward_data,
  input         io_es_dest_valid_es_is_ld,
  input         io_es_dest_valid_es_ready_go,
  input         io_es_dest_valid_es_to_ms_valid,
  input         io_ms_dest_valid_gr_we,
  input         io_ms_dest_valid_ms_valid,
  input  [4:0]  io_ms_dest_valid_dest,
  input  [63:0] io_ms_dest_valid_ms_forward_data,
  input         io_ms_dest_valid_ms_is_ld,
  input         io_ms_dest_valid_ms_to_ws_valid,
  input         io_ms_dest_valid_ms_ready_go,
  input         io_ws_dest_valid_gr_we,
  input         io_ws_dest_valid_ws_valid,
  input  [4:0]  io_ws_dest_valid_dest,
  input  [63:0] io_ws_dest_valid_ws_forward_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  Registers_clock; // @[IDU.scala 283:25]
  wire  Registers_io_wen; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_wdata; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_rdata1; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_rdata2; // @[IDU.scala 283:25]
  wire [4:0] Registers_io_rs1; // @[IDU.scala 283:25]
  wire [4:0] Registers_io_rs2; // @[IDU.scala 283:25]
  wire [4:0] Registers_io_waddr; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_0; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_1; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_2; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_3; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_4; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_5; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_6; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_7; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_8; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_9; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_10; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_11; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_12; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_13; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_14; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_15; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_16; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_17; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_18; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_19; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_20; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_21; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_22; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_23; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_24; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_25; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_26; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_27; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_28; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_29; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_30; // @[IDU.scala 283:25]
  wire [63:0] Registers_io_regs_31; // @[IDU.scala 283:25]
  wire [31:0] DPI_EBREAK_flag; // @[IDU.scala 306:26]
  wire  CSR_clock; // @[IDU.scala 310:20]
  wire  CSR_io_wen; // @[IDU.scala 310:20]
  wire  CSR_io_ren; // @[IDU.scala 310:20]
  wire [63:0] CSR_io_wdata1; // @[IDU.scala 310:20]
  wire [63:0] CSR_io_wdata2; // @[IDU.scala 310:20]
  wire [63:0] CSR_io_rdata; // @[IDU.scala 310:20]
  wire [4:0] CSR_io_waddr1; // @[IDU.scala 310:20]
  wire [4:0] CSR_io_waddr2; // @[IDU.scala 310:20]
  wire [4:0] CSR_io_raddr; // @[IDU.scala 310:20]
  wire [63:0] CSR_io_csrs_0; // @[IDU.scala 310:20]
  wire [63:0] CSR_io_csrs_1; // @[IDU.scala 310:20]
  wire [63:0] CSR_io_csrs_2; // @[IDU.scala 310:20]
  wire [63:0] CSR_io_csrs_3; // @[IDU.scala 310:20]
  wire [63:0] CSR_io_csrs_4; // @[IDU.scala 310:20]
  wire [63:0] dpi_rf_0; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_1; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_2; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_3; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_4; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_5; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_6; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_7; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_8; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_9; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_10; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_11; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_12; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_13; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_14; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_15; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_16; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_17; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_18; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_19; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_20; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_21; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_22; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_23; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_24; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_25; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_26; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_27; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_28; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_29; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_30; // @[IDU.scala 323:19]
  wire [63:0] dpi_rf_31; // @[IDU.scala 323:19]
  wire [63:0] dpi_csr_0; // @[IDU.scala 323:19]
  wire [63:0] dpi_csr_1; // @[IDU.scala 323:19]
  wire [63:0] dpi_csr_2; // @[IDU.scala 323:19]
  wire [63:0] dpi_csr_3; // @[IDU.scala 323:19]
  wire [63:0] dpi_csr_4; // @[IDU.scala 323:19]
  wire [31:0] dpi_inst; // @[IDU.scala 323:19]
  wire [63:0] dpi_pc; // @[IDU.scala 323:19]
  wire [31:0] dpi_eval; // @[IDU.scala 323:19]
  reg  ds_valid; // @[IDU.scala 31:28]
  reg [31:0] fd_bus_r_inst; // @[IDU.scala 33:28]
  reg [31:0] fd_bus_r_pc; // @[IDU.scala 33:28]
  wire [4:0] rs1 = fd_bus_r_inst[19:15]; // @[IDU.scala 269:17]
  wire [4:0] rs2 = fd_bus_r_inst[24:20]; // @[IDU.scala 270:17]
  wire  _es_rawblock_T_1 = rs2 == io_es_dest_valid_dest; // @[IDU.scala 275:59]
  wire  _es_rawblock_T_3 = io_es_dest_valid_dest != 5'h0; // @[IDU.scala 275:111]
  wire  es_rawblock = (rs1 == io_es_dest_valid_dest | rs2 == io_es_dest_valid_dest) & io_es_dest_valid_dest != 5'h0 &
    io_es_dest_valid_es_is_ld & ds_valid; // @[IDU.scala 275:150]
  wire  _ms_rawblock_T_1 = rs2 == io_ms_dest_valid_dest; // @[IDU.scala 276:59]
  wire  _ms_rawblock_T_3 = io_ms_dest_valid_dest != 5'h0; // @[IDU.scala 276:111]
  wire  ms_rawblock = (rs1 == io_ms_dest_valid_dest | rs2 == io_ms_dest_valid_dest) & io_ms_dest_valid_dest != 5'h0 &
    io_ms_dest_valid_ms_is_ld & ds_valid; // @[IDU.scala 276:150]
  wire  rawblock = io_es_dest_valid_es_valid & es_rawblock | io_ms_dest_valid_ms_valid & ms_rawblock; // @[IDU.scala 277:56]
  wire  ds_ready_go = ~rawblock; // @[IDU.scala 278:18]
  wire  _io_ds_to_es_valid_T = ds_valid & ds_ready_go; // @[IDU.scala 56:33]
  wire  eval = io_de_bus_OP == 8'h3f; // @[IDU.scala 226:27]
  wire  mret = io_de_bus_OP == 8'h40; // @[IDU.scala 227:27]
  wire  _br_taken_cancel_T = eval | mret; // @[IDU.scala 267:28]
  wire  _rf_rdata1_T_5 = Registers_io_rs1 == io_es_dest_valid_dest & _es_rawblock_T_3 & io_es_dest_valid_es_to_ms_valid
     & io_es_dest_valid_gr_we & io_es_dest_valid_es_ready_go; // @[IDU.scala 292:144]
  wire  _rf_rdata1_T_11 = Registers_io_rs1 == io_ms_dest_valid_dest & _ms_rawblock_T_3 & io_ms_dest_valid_ms_to_ws_valid
     & io_ms_dest_valid_gr_we & io_ms_dest_valid_ms_ready_go; // @[IDU.scala 293:144]
  wire  _rf_rdata1_T_13 = io_ws_dest_valid_dest != 5'h0; // @[IDU.scala 294:74]
  wire  _rf_rdata1_T_16 = Registers_io_rs1 == io_ws_dest_valid_dest & io_ws_dest_valid_dest != 5'h0 &
    io_ws_dest_valid_ws_valid & io_ws_dest_valid_gr_we; // @[IDU.scala 294:112]
  wire [63:0] _rf_rdata1_T_17 = _rf_rdata1_T_16 ? io_ws_dest_valid_ws_forward_data : Registers_io_rdata1; // @[Mux.scala 101:16]
  wire [63:0] _rf_rdata1_T_18 = _rf_rdata1_T_11 ? io_ms_dest_valid_ms_forward_data : _rf_rdata1_T_17; // @[Mux.scala 101:16]
  wire [63:0] rf_rdata1 = _rf_rdata1_T_5 ? io_es_dest_valid_es_forward_data : _rf_rdata1_T_18; // @[Mux.scala 101:16]
  wire  _rf_rdata2_T_5 = _es_rawblock_T_1 & _es_rawblock_T_3 & io_es_dest_valid_es_to_ms_valid & io_es_dest_valid_gr_we
     & io_es_dest_valid_es_ready_go; // @[IDU.scala 300:136]
  wire  _rf_rdata2_T_11 = _ms_rawblock_T_1 & _ms_rawblock_T_3 & io_ms_dest_valid_ms_to_ws_valid & io_ms_dest_valid_gr_we
     & io_ms_dest_valid_ms_ready_go; // @[IDU.scala 301:134]
  wire  _rf_rdata2_T_16 = rs2 == io_ws_dest_valid_dest & _rf_rdata1_T_13 & io_ws_dest_valid_ws_valid &
    io_ws_dest_valid_gr_we; // @[IDU.scala 302:102]
  wire [63:0] _rf_rdata2_T_17 = _rf_rdata2_T_16 ? io_ws_dest_valid_ws_forward_data : Registers_io_rdata2; // @[Mux.scala 101:16]
  wire [63:0] _rf_rdata2_T_18 = _rf_rdata2_T_11 ? io_ms_dest_valid_ms_forward_data : _rf_rdata2_T_17; // @[Mux.scala 101:16]
  wire [63:0] rf_rdata2 = _rf_rdata2_T_5 ? io_es_dest_valid_es_forward_data : _rf_rdata2_T_18; // @[Mux.scala 101:16]
  wire  _br_taken_T_27 = rf_rdata1 >= rf_rdata2 & ds_valid & ds_ready_go; // @[IDU.scala 247:57]
  wire  _br_taken_T_23 = rf_rdata1 < rf_rdata2 & ds_valid & ds_ready_go; // @[IDU.scala 246:56]
  wire [63:0] _br_taken_T_14 = _rf_rdata1_T_5 ? io_es_dest_valid_es_forward_data : _rf_rdata1_T_18; // @[IDU.scala 245:30]
  wire [63:0] _br_taken_T_15 = _rf_rdata2_T_5 ? io_es_dest_valid_es_forward_data : _rf_rdata2_T_18; // @[IDU.scala 245:50]
  wire  _br_taken_T_19 = $signed(_br_taken_T_14) >= $signed(_br_taken_T_15) & ds_valid & ds_ready_go; // @[IDU.scala 245:70]
  wire  _br_taken_T_13 = $signed(_br_taken_T_14) < $signed(_br_taken_T_15) & ds_valid & ds_ready_go; // @[IDU.scala 244:69]
  wire  _br_taken_T_7 = rf_rdata1 != rf_rdata2 & ds_valid & ds_ready_go; // @[IDU.scala 243:57]
  wire  _br_taken_T_3 = rf_rdata1 == rf_rdata2 & ds_valid & ds_ready_go; // @[IDU.scala 242:57]
  wire  _br_taken_T_37 = 8'h33 == io_de_bus_OP ? _br_taken_T_7 : 8'h32 == io_de_bus_OP & _br_taken_T_3; // @[Mux.scala 81:58]
  wire  _br_taken_T_39 = 8'h36 == io_de_bus_OP ? _br_taken_T_13 : _br_taken_T_37; // @[Mux.scala 81:58]
  wire  _br_taken_T_41 = 8'h34 == io_de_bus_OP ? _br_taken_T_19 : _br_taken_T_39; // @[Mux.scala 81:58]
  wire  _br_taken_T_43 = 8'h37 == io_de_bus_OP ? _br_taken_T_23 : _br_taken_T_41; // @[Mux.scala 81:58]
  wire  _br_taken_T_45 = 8'h35 == io_de_bus_OP ? _br_taken_T_27 : _br_taken_T_43; // @[Mux.scala 81:58]
  wire  _br_taken_T_47 = 8'h3a == io_de_bus_OP ? _io_ds_to_es_valid_T : _br_taken_T_45; // @[Mux.scala 81:58]
  wire  br_taken = 8'h1b == io_de_bus_OP ? _io_ds_to_es_valid_T : _br_taken_T_47; // @[Mux.scala 81:58]
  wire  br_taken_cancel = (eval | mret | br_taken) & ds_ready_go; // @[IDU.scala 267:49]
  wire [31:0] _crtlsignals_T = fd_bus_r_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_1 = 32'h33 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_3 = 32'h3b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_5 = 32'h40000033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_7 = 32'h4000003b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_9 = 32'h2000033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_11 = 32'h200003b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_13 = 32'h2004033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_15 = 32'h2005033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_17 = 32'h200403b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_19 = 32'h200503b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_21 = 32'h1033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_23 = 32'h2033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_25 = 32'h3033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_27 = 32'h103b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_29 = 32'h40005033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_31 = 32'h4000503b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_33 = 32'h5033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_35 = 32'h503b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_37 = 32'h4033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_39 = 32'h7033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_41 = 32'h6033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_43 = 32'h2006033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_45 = 32'h2007033 == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_47 = 32'h200603b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_49 = 32'h200703b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire [31:0] _crtlsignals_T_50 = fd_bus_r_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_51 = 32'h13 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_53 = 32'h1b == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_55 = 32'h67 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_57 = 32'h3 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_59 = 32'h4003 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_61 = 32'h1003 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_63 = 32'h5003 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_65 = 32'h2003 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_67 = 32'h6003 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_69 = 32'h3003 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire [31:0] _crtlsignals_T_70 = fd_bus_r_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_71 = 32'h1013 == _crtlsignals_T_70; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_73 = 32'h101b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_75 = 32'h5013 == _crtlsignals_T_70; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_77 = 32'h501b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_79 = 32'h2013 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_81 = 32'h3013 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_83 = 32'h7013 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_85 = 32'h4013 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_87 = 32'h6013 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_89 = 32'h40005013 == _crtlsignals_T_70; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_91 = 32'h4000501b == _crtlsignals_T; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_93 = 32'h1073 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_95 = 32'h2073 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_97 = 32'h3073 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_99 = 32'h73 == fd_bus_r_inst; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_101 = 32'h3023 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_103 = 32'h23 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_105 = 32'h1023 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_107 = 32'h2023 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_109 = 32'h63 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_111 = 32'h1063 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_113 = 32'h4063 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_115 = 32'h5063 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_117 = 32'h7063 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_119 = 32'h6063 == _crtlsignals_T_50; // @[Lookup.scala 31:38]
  wire [31:0] _crtlsignals_T_120 = fd_bus_r_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_121 = 32'h37 == _crtlsignals_T_120; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_123 = 32'h17 == _crtlsignals_T_120; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_125 = 32'h6f == _crtlsignals_T_120; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_127 = 32'h30200073 == fd_bus_r_inst; // @[Lookup.scala 31:38]
  wire  _crtlsignals_T_129 = 32'h100073 == fd_bus_r_inst; // @[Lookup.scala 31:38]
  wire [7:0] _crtlsignals_T_133 = _crtlsignals_T_129 ? 8'h3b : 8'hff; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_134 = _crtlsignals_T_127 ? 8'h40 : _crtlsignals_T_133; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_135 = _crtlsignals_T_125 ? 8'h3a : _crtlsignals_T_134; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_136 = _crtlsignals_T_123 ? 8'h39 : _crtlsignals_T_135; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_137 = _crtlsignals_T_121 ? 8'h38 : _crtlsignals_T_136; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_138 = _crtlsignals_T_119 ? 8'h37 : _crtlsignals_T_137; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_139 = _crtlsignals_T_117 ? 8'h35 : _crtlsignals_T_138; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_140 = _crtlsignals_T_115 ? 8'h34 : _crtlsignals_T_139; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_141 = _crtlsignals_T_113 ? 8'h36 : _crtlsignals_T_140; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_142 = _crtlsignals_T_111 ? 8'h33 : _crtlsignals_T_141; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_143 = _crtlsignals_T_109 ? 8'h32 : _crtlsignals_T_142; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_144 = _crtlsignals_T_107 ? 8'h31 : _crtlsignals_T_143; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_145 = _crtlsignals_T_105 ? 8'h30 : _crtlsignals_T_144; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_146 = _crtlsignals_T_103 ? 8'h2f : _crtlsignals_T_145; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_147 = _crtlsignals_T_101 ? 8'h2e : _crtlsignals_T_146; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_148 = _crtlsignals_T_99 ? 8'h3f : _crtlsignals_T_147; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_149 = _crtlsignals_T_97 ? 8'h3e : _crtlsignals_T_148; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_150 = _crtlsignals_T_95 ? 8'h3d : _crtlsignals_T_149; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_151 = _crtlsignals_T_93 ? 8'h3c : _crtlsignals_T_150; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_152 = _crtlsignals_T_91 ? 8'h28 : _crtlsignals_T_151; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_153 = _crtlsignals_T_89 ? 8'h27 : _crtlsignals_T_152; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_154 = _crtlsignals_T_87 ? 8'h2d : _crtlsignals_T_153; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_155 = _crtlsignals_T_85 ? 8'h2c : _crtlsignals_T_154; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_156 = _crtlsignals_T_83 ? 8'h2b : _crtlsignals_T_155; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_157 = _crtlsignals_T_81 ? 8'h2a : _crtlsignals_T_156; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_158 = _crtlsignals_T_79 ? 8'h29 : _crtlsignals_T_157; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_159 = _crtlsignals_T_77 ? 8'h26 : _crtlsignals_T_158; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_160 = _crtlsignals_T_75 ? 8'h25 : _crtlsignals_T_159; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_161 = _crtlsignals_T_73 ? 8'h24 : _crtlsignals_T_160; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_162 = _crtlsignals_T_71 ? 8'h23 : _crtlsignals_T_161; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_163 = _crtlsignals_T_69 ? 8'h20 : _crtlsignals_T_162; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_164 = _crtlsignals_T_67 ? 8'h22 : _crtlsignals_T_163; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_165 = _crtlsignals_T_65 ? 8'h21 : _crtlsignals_T_164; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_166 = _crtlsignals_T_63 ? 8'h1f : _crtlsignals_T_165; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_167 = _crtlsignals_T_61 ? 8'h1e : _crtlsignals_T_166; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_168 = _crtlsignals_T_59 ? 8'h1d : _crtlsignals_T_167; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_169 = _crtlsignals_T_57 ? 8'h1c : _crtlsignals_T_168; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_170 = _crtlsignals_T_55 ? 8'h1b : _crtlsignals_T_169; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_171 = _crtlsignals_T_53 ? 8'h1a : _crtlsignals_T_170; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_172 = _crtlsignals_T_51 ? 8'h19 : _crtlsignals_T_171; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_173 = _crtlsignals_T_49 ? 8'h18 : _crtlsignals_T_172; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_174 = _crtlsignals_T_47 ? 8'h17 : _crtlsignals_T_173; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_175 = _crtlsignals_T_45 ? 8'h16 : _crtlsignals_T_174; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_176 = _crtlsignals_T_43 ? 8'h15 : _crtlsignals_T_175; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_177 = _crtlsignals_T_41 ? 8'h14 : _crtlsignals_T_176; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_178 = _crtlsignals_T_39 ? 8'h12 : _crtlsignals_T_177; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_179 = _crtlsignals_T_37 ? 8'h11 : _crtlsignals_T_178; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_180 = _crtlsignals_T_35 ? 8'h10 : _crtlsignals_T_179; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_181 = _crtlsignals_T_33 ? 8'hf : _crtlsignals_T_180; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_182 = _crtlsignals_T_31 ? 8'he : _crtlsignals_T_181; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_183 = _crtlsignals_T_29 ? 8'h13 : _crtlsignals_T_182; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_184 = _crtlsignals_T_27 ? 8'hd : _crtlsignals_T_183; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_185 = _crtlsignals_T_25 ? 8'hc : _crtlsignals_T_184; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_186 = _crtlsignals_T_23 ? 8'hb : _crtlsignals_T_185; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_187 = _crtlsignals_T_21 ? 8'ha : _crtlsignals_T_186; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_188 = _crtlsignals_T_19 ? 8'h9 : _crtlsignals_T_187; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_189 = _crtlsignals_T_17 ? 8'h8 : _crtlsignals_T_188; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_190 = _crtlsignals_T_15 ? 8'h7 : _crtlsignals_T_189; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_191 = _crtlsignals_T_13 ? 8'h6 : _crtlsignals_T_190; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_192 = _crtlsignals_T_11 ? 8'h5 : _crtlsignals_T_191; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_193 = _crtlsignals_T_9 ? 8'h4 : _crtlsignals_T_192; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_194 = _crtlsignals_T_7 ? 8'h3 : _crtlsignals_T_193; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_195 = _crtlsignals_T_5 ? 8'h2 : _crtlsignals_T_194; // @[Lookup.scala 34:39]
  wire [7:0] _crtlsignals_T_196 = _crtlsignals_T_3 ? 8'h1 : _crtlsignals_T_195; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_203 = _crtlsignals_T_119 ? 1'h0 : _crtlsignals_T_121 | (_crtlsignals_T_123 | _crtlsignals_T_125); // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_204 = _crtlsignals_T_117 ? 1'h0 : _crtlsignals_T_203; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_205 = _crtlsignals_T_115 ? 1'h0 : _crtlsignals_T_204; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_206 = _crtlsignals_T_113 ? 1'h0 : _crtlsignals_T_205; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_207 = _crtlsignals_T_111 ? 1'h0 : _crtlsignals_T_206; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_208 = _crtlsignals_T_109 ? 1'h0 : _crtlsignals_T_207; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_209 = _crtlsignals_T_107 ? 1'h0 : _crtlsignals_T_208; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_210 = _crtlsignals_T_105 ? 1'h0 : _crtlsignals_T_209; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_211 = _crtlsignals_T_103 ? 1'h0 : _crtlsignals_T_210; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_212 = _crtlsignals_T_101 ? 1'h0 : _crtlsignals_T_211; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_242 = _crtlsignals_T_41 | (_crtlsignals_T_43 | (_crtlsignals_T_45 | (_crtlsignals_T_47 | (
    _crtlsignals_T_49 | (_crtlsignals_T_51 | (_crtlsignals_T_53 | (_crtlsignals_T_55 | (_crtlsignals_T_57 | (
    _crtlsignals_T_59 | (_crtlsignals_T_61 | (_crtlsignals_T_63 | (_crtlsignals_T_65 | (_crtlsignals_T_67 | (
    _crtlsignals_T_69 | (_crtlsignals_T_71 | (_crtlsignals_T_73 | (_crtlsignals_T_75 | (_crtlsignals_T_77 | (
    _crtlsignals_T_79 | (_crtlsignals_T_81 | (_crtlsignals_T_83 | (_crtlsignals_T_85 | (_crtlsignals_T_87 | (
    _crtlsignals_T_89 | (_crtlsignals_T_91 | (_crtlsignals_T_93 | (_crtlsignals_T_95 | (_crtlsignals_T_97 | (
    _crtlsignals_T_99 | _crtlsignals_T_212))))))))))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_265 = _crtlsignals_T_125 ? 3'h4 : 3'h0; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_266 = _crtlsignals_T_123 ? 3'h3 : _crtlsignals_T_265; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_267 = _crtlsignals_T_121 ? 3'h3 : _crtlsignals_T_266; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_268 = _crtlsignals_T_119 ? 3'h2 : _crtlsignals_T_267; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_269 = _crtlsignals_T_117 ? 3'h2 : _crtlsignals_T_268; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_270 = _crtlsignals_T_115 ? 3'h2 : _crtlsignals_T_269; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_271 = _crtlsignals_T_113 ? 3'h2 : _crtlsignals_T_270; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_272 = _crtlsignals_T_111 ? 3'h2 : _crtlsignals_T_271; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_273 = _crtlsignals_T_109 ? 3'h2 : _crtlsignals_T_272; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_274 = _crtlsignals_T_107 ? 3'h1 : _crtlsignals_T_273; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_275 = _crtlsignals_T_105 ? 3'h1 : _crtlsignals_T_274; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_276 = _crtlsignals_T_103 ? 3'h1 : _crtlsignals_T_275; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_277 = _crtlsignals_T_101 ? 3'h1 : _crtlsignals_T_276; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_278 = _crtlsignals_T_99 ? 3'h0 : _crtlsignals_T_277; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_279 = _crtlsignals_T_97 ? 3'h0 : _crtlsignals_T_278; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_280 = _crtlsignals_T_95 ? 3'h0 : _crtlsignals_T_279; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_281 = _crtlsignals_T_93 ? 3'h0 : _crtlsignals_T_280; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_282 = _crtlsignals_T_91 ? 3'h0 : _crtlsignals_T_281; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_283 = _crtlsignals_T_89 ? 3'h0 : _crtlsignals_T_282; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_284 = _crtlsignals_T_87 ? 3'h0 : _crtlsignals_T_283; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_285 = _crtlsignals_T_85 ? 3'h0 : _crtlsignals_T_284; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_286 = _crtlsignals_T_83 ? 3'h0 : _crtlsignals_T_285; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_287 = _crtlsignals_T_81 ? 3'h0 : _crtlsignals_T_286; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_288 = _crtlsignals_T_79 ? 3'h0 : _crtlsignals_T_287; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_289 = _crtlsignals_T_77 ? 3'h0 : _crtlsignals_T_288; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_290 = _crtlsignals_T_75 ? 3'h0 : _crtlsignals_T_289; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_291 = _crtlsignals_T_73 ? 3'h0 : _crtlsignals_T_290; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_292 = _crtlsignals_T_71 ? 3'h0 : _crtlsignals_T_291; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_293 = _crtlsignals_T_69 ? 3'h0 : _crtlsignals_T_292; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_294 = _crtlsignals_T_67 ? 3'h0 : _crtlsignals_T_293; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_295 = _crtlsignals_T_65 ? 3'h0 : _crtlsignals_T_294; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_296 = _crtlsignals_T_63 ? 3'h0 : _crtlsignals_T_295; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_297 = _crtlsignals_T_61 ? 3'h0 : _crtlsignals_T_296; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_298 = _crtlsignals_T_59 ? 3'h0 : _crtlsignals_T_297; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_299 = _crtlsignals_T_57 ? 3'h0 : _crtlsignals_T_298; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_300 = _crtlsignals_T_55 ? 3'h0 : _crtlsignals_T_299; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_301 = _crtlsignals_T_53 ? 3'h0 : _crtlsignals_T_300; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_302 = _crtlsignals_T_51 ? 3'h0 : _crtlsignals_T_301; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_303 = _crtlsignals_T_49 ? 3'h0 : _crtlsignals_T_302; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_304 = _crtlsignals_T_47 ? 3'h0 : _crtlsignals_T_303; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_305 = _crtlsignals_T_45 ? 3'h0 : _crtlsignals_T_304; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_306 = _crtlsignals_T_43 ? 3'h0 : _crtlsignals_T_305; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_307 = _crtlsignals_T_41 ? 3'h0 : _crtlsignals_T_306; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_308 = _crtlsignals_T_39 ? 3'h0 : _crtlsignals_T_307; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_309 = _crtlsignals_T_37 ? 3'h0 : _crtlsignals_T_308; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_310 = _crtlsignals_T_35 ? 3'h0 : _crtlsignals_T_309; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_311 = _crtlsignals_T_33 ? 3'h0 : _crtlsignals_T_310; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_312 = _crtlsignals_T_31 ? 3'h0 : _crtlsignals_T_311; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_313 = _crtlsignals_T_29 ? 3'h0 : _crtlsignals_T_312; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_314 = _crtlsignals_T_27 ? 3'h0 : _crtlsignals_T_313; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_315 = _crtlsignals_T_25 ? 3'h0 : _crtlsignals_T_314; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_316 = _crtlsignals_T_23 ? 3'h0 : _crtlsignals_T_315; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_317 = _crtlsignals_T_21 ? 3'h0 : _crtlsignals_T_316; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_318 = _crtlsignals_T_19 ? 3'h0 : _crtlsignals_T_317; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_319 = _crtlsignals_T_17 ? 3'h0 : _crtlsignals_T_318; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_320 = _crtlsignals_T_15 ? 3'h0 : _crtlsignals_T_319; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_321 = _crtlsignals_T_13 ? 3'h0 : _crtlsignals_T_320; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_322 = _crtlsignals_T_11 ? 3'h0 : _crtlsignals_T_321; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_323 = _crtlsignals_T_9 ? 3'h0 : _crtlsignals_T_322; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_324 = _crtlsignals_T_7 ? 3'h0 : _crtlsignals_T_323; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_325 = _crtlsignals_T_5 ? 3'h0 : _crtlsignals_T_324; // @[Lookup.scala 34:39]
  wire [2:0] _crtlsignals_T_326 = _crtlsignals_T_3 ? 3'h0 : _crtlsignals_T_325; // @[Lookup.scala 34:39]
  wire [2:0] ImmType = _crtlsignals_T_1 ? 3'h0 : _crtlsignals_T_326; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_408 = _crtlsignals_T_99 ? 1'h0 : _crtlsignals_T_101 | (_crtlsignals_T_103 | (_crtlsignals_T_105
     | _crtlsignals_T_107)); // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_409 = _crtlsignals_T_97 ? 1'h0 : _crtlsignals_T_408; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_410 = _crtlsignals_T_95 ? 1'h0 : _crtlsignals_T_409; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_411 = _crtlsignals_T_93 ? 1'h0 : _crtlsignals_T_410; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_412 = _crtlsignals_T_91 ? 1'h0 : _crtlsignals_T_411; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_413 = _crtlsignals_T_89 ? 1'h0 : _crtlsignals_T_412; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_414 = _crtlsignals_T_87 ? 1'h0 : _crtlsignals_T_413; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_415 = _crtlsignals_T_85 ? 1'h0 : _crtlsignals_T_414; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_416 = _crtlsignals_T_83 ? 1'h0 : _crtlsignals_T_415; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_417 = _crtlsignals_T_81 ? 1'h0 : _crtlsignals_T_416; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_418 = _crtlsignals_T_79 ? 1'h0 : _crtlsignals_T_417; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_419 = _crtlsignals_T_77 ? 1'h0 : _crtlsignals_T_418; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_420 = _crtlsignals_T_75 ? 1'h0 : _crtlsignals_T_419; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_421 = _crtlsignals_T_73 ? 1'h0 : _crtlsignals_T_420; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_422 = _crtlsignals_T_71 ? 1'h0 : _crtlsignals_T_421; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_423 = _crtlsignals_T_69 ? 1'h0 : _crtlsignals_T_422; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_424 = _crtlsignals_T_67 ? 1'h0 : _crtlsignals_T_423; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_425 = _crtlsignals_T_65 ? 1'h0 : _crtlsignals_T_424; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_426 = _crtlsignals_T_63 ? 1'h0 : _crtlsignals_T_425; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_427 = _crtlsignals_T_61 ? 1'h0 : _crtlsignals_T_426; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_428 = _crtlsignals_T_59 ? 1'h0 : _crtlsignals_T_427; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_429 = _crtlsignals_T_57 ? 1'h0 : _crtlsignals_T_428; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_430 = _crtlsignals_T_55 ? 1'h0 : _crtlsignals_T_429; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_431 = _crtlsignals_T_53 ? 1'h0 : _crtlsignals_T_430; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_432 = _crtlsignals_T_51 ? 1'h0 : _crtlsignals_T_431; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_433 = _crtlsignals_T_49 ? 1'h0 : _crtlsignals_T_432; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_434 = _crtlsignals_T_47 ? 1'h0 : _crtlsignals_T_433; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_435 = _crtlsignals_T_45 ? 1'h0 : _crtlsignals_T_434; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_436 = _crtlsignals_T_43 ? 1'h0 : _crtlsignals_T_435; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_437 = _crtlsignals_T_41 ? 1'h0 : _crtlsignals_T_436; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_438 = _crtlsignals_T_39 ? 1'h0 : _crtlsignals_T_437; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_439 = _crtlsignals_T_37 ? 1'h0 : _crtlsignals_T_438; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_440 = _crtlsignals_T_35 ? 1'h0 : _crtlsignals_T_439; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_441 = _crtlsignals_T_33 ? 1'h0 : _crtlsignals_T_440; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_442 = _crtlsignals_T_31 ? 1'h0 : _crtlsignals_T_441; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_443 = _crtlsignals_T_29 ? 1'h0 : _crtlsignals_T_442; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_444 = _crtlsignals_T_27 ? 1'h0 : _crtlsignals_T_443; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_445 = _crtlsignals_T_25 ? 1'h0 : _crtlsignals_T_444; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_446 = _crtlsignals_T_23 ? 1'h0 : _crtlsignals_T_445; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_447 = _crtlsignals_T_21 ? 1'h0 : _crtlsignals_T_446; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_448 = _crtlsignals_T_19 ? 1'h0 : _crtlsignals_T_447; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_449 = _crtlsignals_T_17 ? 1'h0 : _crtlsignals_T_448; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_450 = _crtlsignals_T_15 ? 1'h0 : _crtlsignals_T_449; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_451 = _crtlsignals_T_13 ? 1'h0 : _crtlsignals_T_450; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_452 = _crtlsignals_T_11 ? 1'h0 : _crtlsignals_T_451; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_453 = _crtlsignals_T_9 ? 1'h0 : _crtlsignals_T_452; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_454 = _crtlsignals_T_7 ? 1'h0 : _crtlsignals_T_453; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_455 = _crtlsignals_T_5 ? 1'h0 : _crtlsignals_T_454; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_456 = _crtlsignals_T_3 ? 1'h0 : _crtlsignals_T_455; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_495 = _crtlsignals_T_55 ? 1'h0 : _crtlsignals_T_57 | (_crtlsignals_T_59 | (_crtlsignals_T_61 | (
    _crtlsignals_T_63 | (_crtlsignals_T_65 | (_crtlsignals_T_67 | _crtlsignals_T_69))))); // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_496 = _crtlsignals_T_53 ? 1'h0 : _crtlsignals_T_495; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_497 = _crtlsignals_T_51 ? 1'h0 : _crtlsignals_T_496; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_498 = _crtlsignals_T_49 ? 1'h0 : _crtlsignals_T_497; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_499 = _crtlsignals_T_47 ? 1'h0 : _crtlsignals_T_498; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_500 = _crtlsignals_T_45 ? 1'h0 : _crtlsignals_T_499; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_501 = _crtlsignals_T_43 ? 1'h0 : _crtlsignals_T_500; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_502 = _crtlsignals_T_41 ? 1'h0 : _crtlsignals_T_501; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_503 = _crtlsignals_T_39 ? 1'h0 : _crtlsignals_T_502; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_504 = _crtlsignals_T_37 ? 1'h0 : _crtlsignals_T_503; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_505 = _crtlsignals_T_35 ? 1'h0 : _crtlsignals_T_504; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_506 = _crtlsignals_T_33 ? 1'h0 : _crtlsignals_T_505; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_507 = _crtlsignals_T_31 ? 1'h0 : _crtlsignals_T_506; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_508 = _crtlsignals_T_29 ? 1'h0 : _crtlsignals_T_507; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_509 = _crtlsignals_T_27 ? 1'h0 : _crtlsignals_T_508; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_510 = _crtlsignals_T_25 ? 1'h0 : _crtlsignals_T_509; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_511 = _crtlsignals_T_23 ? 1'h0 : _crtlsignals_T_510; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_512 = _crtlsignals_T_21 ? 1'h0 : _crtlsignals_T_511; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_513 = _crtlsignals_T_19 ? 1'h0 : _crtlsignals_T_512; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_514 = _crtlsignals_T_17 ? 1'h0 : _crtlsignals_T_513; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_515 = _crtlsignals_T_15 ? 1'h0 : _crtlsignals_T_514; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_516 = _crtlsignals_T_13 ? 1'h0 : _crtlsignals_T_515; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_517 = _crtlsignals_T_11 ? 1'h0 : _crtlsignals_T_516; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_518 = _crtlsignals_T_9 ? 1'h0 : _crtlsignals_T_517; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_519 = _crtlsignals_T_7 ? 1'h0 : _crtlsignals_T_518; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_520 = _crtlsignals_T_5 ? 1'h0 : _crtlsignals_T_519; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_521 = _crtlsignals_T_3 ? 1'h0 : _crtlsignals_T_520; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_542 = _crtlsignals_T_91 ? 1'h0 : _crtlsignals_T_93 | (_crtlsignals_T_95 | (_crtlsignals_T_97 |
    _crtlsignals_T_99)); // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_543 = _crtlsignals_T_89 ? 1'h0 : _crtlsignals_T_542; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_544 = _crtlsignals_T_87 ? 1'h0 : _crtlsignals_T_543; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_545 = _crtlsignals_T_85 ? 1'h0 : _crtlsignals_T_544; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_546 = _crtlsignals_T_83 ? 1'h0 : _crtlsignals_T_545; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_547 = _crtlsignals_T_81 ? 1'h0 : _crtlsignals_T_546; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_548 = _crtlsignals_T_79 ? 1'h0 : _crtlsignals_T_547; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_549 = _crtlsignals_T_77 ? 1'h0 : _crtlsignals_T_548; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_550 = _crtlsignals_T_75 ? 1'h0 : _crtlsignals_T_549; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_551 = _crtlsignals_T_73 ? 1'h0 : _crtlsignals_T_550; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_552 = _crtlsignals_T_71 ? 1'h0 : _crtlsignals_T_551; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_553 = _crtlsignals_T_69 ? 1'h0 : _crtlsignals_T_552; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_554 = _crtlsignals_T_67 ? 1'h0 : _crtlsignals_T_553; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_555 = _crtlsignals_T_65 ? 1'h0 : _crtlsignals_T_554; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_556 = _crtlsignals_T_63 ? 1'h0 : _crtlsignals_T_555; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_557 = _crtlsignals_T_61 ? 1'h0 : _crtlsignals_T_556; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_558 = _crtlsignals_T_59 ? 1'h0 : _crtlsignals_T_557; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_559 = _crtlsignals_T_57 ? 1'h0 : _crtlsignals_T_558; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_560 = _crtlsignals_T_55 ? 1'h0 : _crtlsignals_T_559; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_561 = _crtlsignals_T_53 ? 1'h0 : _crtlsignals_T_560; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_562 = _crtlsignals_T_51 ? 1'h0 : _crtlsignals_T_561; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_563 = _crtlsignals_T_49 ? 1'h0 : _crtlsignals_T_562; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_564 = _crtlsignals_T_47 ? 1'h0 : _crtlsignals_T_563; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_565 = _crtlsignals_T_45 ? 1'h0 : _crtlsignals_T_564; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_566 = _crtlsignals_T_43 ? 1'h0 : _crtlsignals_T_565; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_567 = _crtlsignals_T_41 ? 1'h0 : _crtlsignals_T_566; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_568 = _crtlsignals_T_39 ? 1'h0 : _crtlsignals_T_567; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_569 = _crtlsignals_T_37 ? 1'h0 : _crtlsignals_T_568; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_570 = _crtlsignals_T_35 ? 1'h0 : _crtlsignals_T_569; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_571 = _crtlsignals_T_33 ? 1'h0 : _crtlsignals_T_570; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_572 = _crtlsignals_T_31 ? 1'h0 : _crtlsignals_T_571; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_573 = _crtlsignals_T_29 ? 1'h0 : _crtlsignals_T_572; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_574 = _crtlsignals_T_27 ? 1'h0 : _crtlsignals_T_573; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_575 = _crtlsignals_T_25 ? 1'h0 : _crtlsignals_T_574; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_576 = _crtlsignals_T_23 ? 1'h0 : _crtlsignals_T_575; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_577 = _crtlsignals_T_21 ? 1'h0 : _crtlsignals_T_576; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_578 = _crtlsignals_T_19 ? 1'h0 : _crtlsignals_T_577; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_579 = _crtlsignals_T_17 ? 1'h0 : _crtlsignals_T_578; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_580 = _crtlsignals_T_15 ? 1'h0 : _crtlsignals_T_579; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_581 = _crtlsignals_T_13 ? 1'h0 : _crtlsignals_T_580; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_582 = _crtlsignals_T_11 ? 1'h0 : _crtlsignals_T_581; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_583 = _crtlsignals_T_9 ? 1'h0 : _crtlsignals_T_582; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_584 = _crtlsignals_T_7 ? 1'h0 : _crtlsignals_T_583; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_585 = _crtlsignals_T_5 ? 1'h0 : _crtlsignals_T_584; // @[Lookup.scala 34:39]
  wire  _crtlsignals_T_586 = _crtlsignals_T_3 ? 1'h0 : _crtlsignals_T_585; // @[Lookup.scala 34:39]
  wire [51:0] _I_T_3 = fd_bus_r_inst[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 74:12]
  wire [63:0] I = {_I_T_3,fd_bus_r_inst[31:20]}; // @[Cat.scala 31:58]
  wire [43:0] _U_T_3 = fd_bus_r_inst[31] ? 44'hfffffffffff : 44'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _U_T_4 = {_U_T_3,fd_bus_r_inst[31:12]}; // @[Cat.scala 31:58]
  wire [75:0] U = {_U_T_4, 12'h0}; // @[IDU.scala 177:37]
  wire [56:0] _S_T_3 = fd_bus_r_inst[31] ? 57'h1ffffffffffffff : 57'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _S_T_4 = {_S_T_3,fd_bus_r_inst[31:25]}; // @[Cat.scala 31:58]
  wire [68:0] _S_T_5 = {_S_T_4, 5'h0}; // @[IDU.scala 178:36]
  wire [68:0] _GEN_4 = {{64'd0}, fd_bus_r_inst[11:7]}; // @[IDU.scala 178:41]
  wire [68:0] S = _S_T_5 | _GEN_4; // @[IDU.scala 178:41]
  wire [62:0] _J_T_3 = fd_bus_r_inst[31] ? 63'h7fffffffffffffff : 63'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _J_T_4 = {_J_T_3,fd_bus_r_inst[31]}; // @[Cat.scala 31:58]
  wire [83:0] _J_T_5 = {_J_T_4, 20'h0}; // @[IDU.scala 179:32]
  wire [11:0] _J_T_7 = {fd_bus_r_inst[20], 11'h0}; // @[IDU.scala 179:52]
  wire [83:0] _GEN_5 = {{72'd0}, _J_T_7}; // @[IDU.scala 179:38]
  wire [83:0] _J_T_8 = _J_T_5 | _GEN_5; // @[IDU.scala 179:38]
  wire [19:0] _J_T_10 = {fd_bus_r_inst[19:12], 12'h0}; // @[IDU.scala 179:76]
  wire [83:0] _GEN_6 = {{64'd0}, _J_T_10}; // @[IDU.scala 179:58]
  wire [83:0] _J_T_11 = _J_T_8 | _GEN_6; // @[IDU.scala 179:58]
  wire [10:0] _J_T_13 = {fd_bus_r_inst[30:21], 1'h0}; // @[IDU.scala 179:100]
  wire [83:0] _GEN_7 = {{73'd0}, _J_T_13}; // @[IDU.scala 179:82]
  wire [83:0] J = _J_T_11 | _GEN_7; // @[IDU.scala 179:82]
  wire [75:0] _B_T_5 = {_J_T_4, 12'h0}; // @[IDU.scala 180:32]
  wire [11:0] _B_T_7 = {fd_bus_r_inst[7], 11'h0}; // @[IDU.scala 180:51]
  wire [75:0] _GEN_8 = {{64'd0}, _B_T_7}; // @[IDU.scala 180:38]
  wire [75:0] _B_T_8 = _B_T_5 | _GEN_8; // @[IDU.scala 180:38]
  wire [10:0] _B_T_10 = {fd_bus_r_inst[30:25], 5'h0}; // @[IDU.scala 180:75]
  wire [75:0] _GEN_9 = {{65'd0}, _B_T_10}; // @[IDU.scala 180:57]
  wire [75:0] _B_T_11 = _B_T_8 | _GEN_9; // @[IDU.scala 180:57]
  wire [4:0] _B_T_13 = {fd_bus_r_inst[11:8], 1'h0}; // @[IDU.scala 180:97]
  wire [75:0] _GEN_10 = {{71'd0}, _B_T_13}; // @[IDU.scala 180:80]
  wire [75:0] B = _B_T_11 | _GEN_10; // @[IDU.scala 180:80]
  wire [63:0] _io_de_bus_imm_T_1 = 3'h0 == ImmType ? I : 64'h0; // @[Mux.scala 81:58]
  wire [68:0] _io_de_bus_imm_T_3 = 3'h1 == ImmType ? S : {{5'd0}, _io_de_bus_imm_T_1}; // @[Mux.scala 81:58]
  wire [75:0] _io_de_bus_imm_T_5 = 3'h2 == ImmType ? B : {{7'd0}, _io_de_bus_imm_T_3}; // @[Mux.scala 81:58]
  wire [75:0] _io_de_bus_imm_T_7 = 3'h3 == ImmType ? U : _io_de_bus_imm_T_5; // @[Mux.scala 81:58]
  wire [83:0] _io_de_bus_imm_T_9 = 3'h4 == ImmType ? J : {{8'd0}, _io_de_bus_imm_T_7}; // @[Mux.scala 81:58]
  wire [63:0] _io_de_bus_wmask_T_1 = 8'h2f == io_de_bus_OP ? 64'h1 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _io_de_bus_wmask_T_3 = 8'h30 == io_de_bus_OP ? 64'h3 : _io_de_bus_wmask_T_1; // @[Mux.scala 81:58]
  wire [63:0] _io_de_bus_wmask_T_5 = 8'h31 == io_de_bus_OP ? 64'hf : _io_de_bus_wmask_T_3; // @[Mux.scala 81:58]
  wire [63:0] _io_de_bus_wmask_T_7 = 8'h2e == io_de_bus_OP ? 64'hff : _io_de_bus_wmask_T_5; // @[Mux.scala 81:58]
  wire [2:0] _io_de_bus_ld_type_T_3 = 8'h1e == io_de_bus_OP ? 3'h1 : 3'h0; // @[Mux.scala 81:58]
  wire [2:0] _io_de_bus_ld_type_T_5 = 8'h21 == io_de_bus_OP ? 3'h2 : _io_de_bus_ld_type_T_3; // @[Mux.scala 81:58]
  wire [2:0] _io_de_bus_ld_type_T_7 = 8'h20 == io_de_bus_OP ? 3'h3 : _io_de_bus_ld_type_T_5; // @[Mux.scala 81:58]
  wire [2:0] _io_de_bus_ld_type_T_9 = 8'h1d == io_de_bus_OP ? 3'h4 : _io_de_bus_ld_type_T_7; // @[Mux.scala 81:58]
  wire [2:0] _io_de_bus_ld_type_T_11 = 8'h1f == io_de_bus_OP ? 3'h5 : _io_de_bus_ld_type_T_9; // @[Mux.scala 81:58]
  wire [1:0] _csr_index_T_3 = 64'h341 == I ? 2'h2 : {{1'd0}, 64'h342 == I}; // @[Mux.scala 81:58]
  wire [1:0] _csr_index_T_5 = 64'h300 == I ? 2'h3 : _csr_index_T_3; // @[Mux.scala 81:58]
  wire [2:0] csr_index = 64'h305 == I ? 3'h4 : {{1'd0}, _csr_index_T_5}; // @[Mux.scala 81:58]
  wire [2:0] _io_de_bus_csr_raddr_T = mret ? 3'h2 : csr_index; // @[IDU.scala 229:42]
  wire [63:0] _GEN_11 = {{32'd0}, fd_bus_r_pc}; // @[IDU.scala 256:25]
  wire [63:0] _br_target_T_1 = _GEN_11 + io_de_bus_imm; // @[IDU.scala 256:25]
  wire [63:0] _br_target_T_15 = rf_rdata1 + io_de_bus_imm; // @[IDU.scala 263:31]
  wire [63:0] _br_target_T_16 = _br_target_T_15 & 64'hfffffffffffffffe; // @[IDU.scala 263:48]
  wire [63:0] _br_target_T_18 = 8'h32 == io_de_bus_OP ? _br_target_T_1 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _br_target_T_20 = 8'h33 == io_de_bus_OP ? _br_target_T_1 : _br_target_T_18; // @[Mux.scala 81:58]
  wire [63:0] _br_target_T_22 = 8'h36 == io_de_bus_OP ? _br_target_T_1 : _br_target_T_20; // @[Mux.scala 81:58]
  wire [63:0] _br_target_T_24 = 8'h34 == io_de_bus_OP ? _br_target_T_1 : _br_target_T_22; // @[Mux.scala 81:58]
  wire [63:0] _br_target_T_26 = 8'h37 == io_de_bus_OP ? _br_target_T_1 : _br_target_T_24; // @[Mux.scala 81:58]
  wire [63:0] _br_target_T_28 = 8'h35 == io_de_bus_OP ? _br_target_T_1 : _br_target_T_26; // @[Mux.scala 81:58]
  wire [63:0] _br_target_T_30 = 8'h3a == io_de_bus_OP ? _br_target_T_1 : _br_target_T_28; // @[Mux.scala 81:58]
  wire [63:0] _br_target_T_32 = 8'h1b == io_de_bus_OP ? _br_target_T_16 : _br_target_T_30; // @[Mux.scala 81:58]
  wire [2:0] _T_7 = io_rf_bus_eval ? io_rf_bus_csr_waddr2 : 3'h0; // @[IDU.scala 312:20]
  Registers Registers ( // @[IDU.scala 283:25]
    .clock(Registers_clock),
    .io_wen(Registers_io_wen),
    .io_wdata(Registers_io_wdata),
    .io_rdata1(Registers_io_rdata1),
    .io_rdata2(Registers_io_rdata2),
    .io_rs1(Registers_io_rs1),
    .io_rs2(Registers_io_rs2),
    .io_waddr(Registers_io_waddr),
    .io_regs_0(Registers_io_regs_0),
    .io_regs_1(Registers_io_regs_1),
    .io_regs_2(Registers_io_regs_2),
    .io_regs_3(Registers_io_regs_3),
    .io_regs_4(Registers_io_regs_4),
    .io_regs_5(Registers_io_regs_5),
    .io_regs_6(Registers_io_regs_6),
    .io_regs_7(Registers_io_regs_7),
    .io_regs_8(Registers_io_regs_8),
    .io_regs_9(Registers_io_regs_9),
    .io_regs_10(Registers_io_regs_10),
    .io_regs_11(Registers_io_regs_11),
    .io_regs_12(Registers_io_regs_12),
    .io_regs_13(Registers_io_regs_13),
    .io_regs_14(Registers_io_regs_14),
    .io_regs_15(Registers_io_regs_15),
    .io_regs_16(Registers_io_regs_16),
    .io_regs_17(Registers_io_regs_17),
    .io_regs_18(Registers_io_regs_18),
    .io_regs_19(Registers_io_regs_19),
    .io_regs_20(Registers_io_regs_20),
    .io_regs_21(Registers_io_regs_21),
    .io_regs_22(Registers_io_regs_22),
    .io_regs_23(Registers_io_regs_23),
    .io_regs_24(Registers_io_regs_24),
    .io_regs_25(Registers_io_regs_25),
    .io_regs_26(Registers_io_regs_26),
    .io_regs_27(Registers_io_regs_27),
    .io_regs_28(Registers_io_regs_28),
    .io_regs_29(Registers_io_regs_29),
    .io_regs_30(Registers_io_regs_30),
    .io_regs_31(Registers_io_regs_31)
  );
  DPI_EBREAK DPI_EBREAK ( // @[IDU.scala 306:26]
    .flag(DPI_EBREAK_flag)
  );
  CSR CSR ( // @[IDU.scala 310:20]
    .clock(CSR_clock),
    .io_wen(CSR_io_wen),
    .io_ren(CSR_io_ren),
    .io_wdata1(CSR_io_wdata1),
    .io_wdata2(CSR_io_wdata2),
    .io_rdata(CSR_io_rdata),
    .io_waddr1(CSR_io_waddr1),
    .io_waddr2(CSR_io_waddr2),
    .io_raddr(CSR_io_raddr),
    .io_csrs_0(CSR_io_csrs_0),
    .io_csrs_1(CSR_io_csrs_1),
    .io_csrs_2(CSR_io_csrs_2),
    .io_csrs_3(CSR_io_csrs_3),
    .io_csrs_4(CSR_io_csrs_4)
  );
  DPI dpi ( // @[IDU.scala 323:19]
    .rf_0(dpi_rf_0),
    .rf_1(dpi_rf_1),
    .rf_2(dpi_rf_2),
    .rf_3(dpi_rf_3),
    .rf_4(dpi_rf_4),
    .rf_5(dpi_rf_5),
    .rf_6(dpi_rf_6),
    .rf_7(dpi_rf_7),
    .rf_8(dpi_rf_8),
    .rf_9(dpi_rf_9),
    .rf_10(dpi_rf_10),
    .rf_11(dpi_rf_11),
    .rf_12(dpi_rf_12),
    .rf_13(dpi_rf_13),
    .rf_14(dpi_rf_14),
    .rf_15(dpi_rf_15),
    .rf_16(dpi_rf_16),
    .rf_17(dpi_rf_17),
    .rf_18(dpi_rf_18),
    .rf_19(dpi_rf_19),
    .rf_20(dpi_rf_20),
    .rf_21(dpi_rf_21),
    .rf_22(dpi_rf_22),
    .rf_23(dpi_rf_23),
    .rf_24(dpi_rf_24),
    .rf_25(dpi_rf_25),
    .rf_26(dpi_rf_26),
    .rf_27(dpi_rf_27),
    .rf_28(dpi_rf_28),
    .rf_29(dpi_rf_29),
    .rf_30(dpi_rf_30),
    .rf_31(dpi_rf_31),
    .csr_0(dpi_csr_0),
    .csr_1(dpi_csr_1),
    .csr_2(dpi_csr_2),
    .csr_3(dpi_csr_3),
    .csr_4(dpi_csr_4),
    .inst(dpi_inst),
    .pc(dpi_pc),
    .eval(dpi_eval)
  );
  assign io_ds_allowin = (~ds_valid | ds_ready_go & io_es_allowin) & ds_ready_go; // @[IDU.scala 55:68]
  assign io_ds_to_es_valid = ds_valid & ds_ready_go; // @[IDU.scala 56:33]
  assign io_de_bus_OP = _crtlsignals_T_1 ? 8'h0 : _crtlsignals_T_196; // @[Lookup.scala 34:39]
  assign io_de_bus_res_from_mem = _crtlsignals_T_1 ? 1'h0 : _crtlsignals_T_521; // @[Lookup.scala 34:39]
  assign io_de_bus_gr_we = _crtlsignals_T_1 | (_crtlsignals_T_3 | (_crtlsignals_T_5 | (_crtlsignals_T_7 | (
    _crtlsignals_T_9 | (_crtlsignals_T_11 | (_crtlsignals_T_13 | (_crtlsignals_T_15 | (_crtlsignals_T_17 | (
    _crtlsignals_T_19 | (_crtlsignals_T_21 | (_crtlsignals_T_23 | (_crtlsignals_T_25 | (_crtlsignals_T_27 | (
    _crtlsignals_T_29 | (_crtlsignals_T_31 | (_crtlsignals_T_33 | (_crtlsignals_T_35 | (_crtlsignals_T_37 | (
    _crtlsignals_T_39 | _crtlsignals_T_242))))))))))))))))))); // @[Lookup.scala 34:39]
  assign io_de_bus_MemWen = _crtlsignals_T_1 ? 1'h0 : _crtlsignals_T_456; // @[Lookup.scala 34:39]
  assign io_de_bus_wmask = _io_de_bus_wmask_T_7[7:0]; // @[IDU.scala 193:19]
  assign io_de_bus_ds_pc = fd_bus_r_pc; // @[IDU.scala 36:21 38:11]
  assign io_de_bus_dest = fd_bus_r_inst[11:7]; // @[IDU.scala 271:17]
  assign io_de_bus_imm = _io_de_bus_imm_T_9[63:0]; // @[IDU.scala 182:17]
  assign io_de_bus_rdata1 = _rf_rdata1_T_5 ? io_es_dest_valid_es_forward_data : _rf_rdata1_T_18; // @[Mux.scala 101:16]
  assign io_de_bus_rdata2 = _rf_rdata2_T_5 ? io_es_dest_valid_es_forward_data : _rf_rdata2_T_18; // @[Mux.scala 101:16]
  assign io_de_bus_ld_type = 8'h22 == io_de_bus_OP ? 3'h6 : _io_de_bus_ld_type_T_11; // @[Mux.scala 81:58]
  assign io_de_bus_inst = fd_bus_r_inst; // @[IDU.scala 35:21 37:11]
  assign io_de_bus_csr_rdata = CSR_io_rdata; // @[IDU.scala 318:23]
  assign io_de_bus_csr_waddr1 = eval ? 3'h1 : csr_index; // @[IDU.scala 230:30]
  assign io_de_bus_csr_waddr2 = eval ? 3'h2 : csr_index; // @[IDU.scala 231:30]
  assign io_de_bus_csr_raddr = eval ? 3'h4 : _io_de_bus_csr_raddr_T; // @[IDU.scala 229:29]
  assign io_de_bus_csr_ren = _br_taken_cancel_T | csr_index != 3'h0; // @[IDU.scala 232:40]
  assign io_de_bus_csr_wen = _crtlsignals_T_1 ? 1'h0 : _crtlsignals_T_586; // @[Lookup.scala 34:39]
  assign io_de_bus_eval = io_de_bus_OP == 8'h3f; // @[IDU.scala 226:27]
  assign io_de_bus_is_ld = io_de_bus_res_from_mem; // @[IDU.scala 273:25]
  assign io_br_bus_br_taken = 8'h1b == io_de_bus_OP ? _io_ds_to_es_valid_T : _br_taken_T_47; // @[Mux.scala 81:58]
  assign io_br_bus_br_target = _br_target_T_32[31:0]; // @[IDU.scala 252:13 48:29]
  assign io_br_bus_rawblock = io_es_dest_valid_es_valid & es_rawblock | io_ms_dest_valid_ms_valid & ms_rawblock; // @[IDU.scala 277:56]
  assign io_br_bus_csr_rdata = CSR_io_rdata; // @[IDU.scala 319:23]
  assign io_br_bus_eval = io_de_bus_OP == 8'h3f; // @[IDU.scala 226:27]
  assign io_br_bus_mret = io_de_bus_OP == 8'h40; // @[IDU.scala 227:27]
  assign Registers_clock = clock;
  assign Registers_io_wen = io_rf_bus_rf_we; // @[IDU.scala 40:22 43:12]
  assign Registers_io_wdata = io_rf_bus_rf_wdata; // @[IDU.scala 42:22 45:12]
  assign Registers_io_rs1 = ~eval ? rs1 : 5'h11; // @[IDU.scala 287:25]
  assign Registers_io_rs2 = fd_bus_r_inst[24:20]; // @[IDU.scala 270:17]
  assign Registers_io_waddr = io_rf_bus_rf_waddr; // @[IDU.scala 41:22 44:12]
  assign DPI_EBREAK_flag = io_de_bus_OP == 8'h3b & ds_valid ? 32'h1 : 32'h0; // @[IDU.scala 307:25]
  assign CSR_clock = clock;
  assign CSR_io_wen = io_rf_bus_csr_wen; // @[IDU.scala 317:14]
  assign CSR_io_ren = io_de_bus_csr_ren; // @[IDU.scala 315:14]
  assign CSR_io_wdata1 = io_rf_bus_csr_wdata; // @[IDU.scala 313:15]
  assign CSR_io_wdata2 = {{32'd0}, io_rf_bus_wb_pc}; // @[IDU.scala 314:15]
  assign CSR_io_waddr1 = {{2'd0}, io_rf_bus_csr_waddr1}; // @[IDU.scala 311:14]
  assign CSR_io_waddr2 = {{2'd0}, _T_7}; // @[IDU.scala 312:14]
  assign CSR_io_raddr = {{2'd0}, io_de_bus_csr_raddr}; // @[IDU.scala 316:14]
  assign dpi_rf_0 = Registers_io_regs_0; // @[IDU.scala 324:16]
  assign dpi_rf_1 = Registers_io_regs_1; // @[IDU.scala 325:16]
  assign dpi_rf_2 = Registers_io_regs_2; // @[IDU.scala 326:16]
  assign dpi_rf_3 = Registers_io_regs_3; // @[IDU.scala 327:16]
  assign dpi_rf_4 = Registers_io_regs_4; // @[IDU.scala 328:16]
  assign dpi_rf_5 = Registers_io_regs_5; // @[IDU.scala 329:16]
  assign dpi_rf_6 = Registers_io_regs_6; // @[IDU.scala 330:16]
  assign dpi_rf_7 = Registers_io_regs_7; // @[IDU.scala 331:16]
  assign dpi_rf_8 = Registers_io_regs_8; // @[IDU.scala 332:16]
  assign dpi_rf_9 = Registers_io_regs_9; // @[IDU.scala 333:16]
  assign dpi_rf_10 = Registers_io_regs_10; // @[IDU.scala 334:16]
  assign dpi_rf_11 = Registers_io_regs_11; // @[IDU.scala 335:16]
  assign dpi_rf_12 = Registers_io_regs_12; // @[IDU.scala 336:16]
  assign dpi_rf_13 = Registers_io_regs_13; // @[IDU.scala 337:16]
  assign dpi_rf_14 = Registers_io_regs_14; // @[IDU.scala 338:16]
  assign dpi_rf_15 = Registers_io_regs_15; // @[IDU.scala 339:16]
  assign dpi_rf_16 = Registers_io_regs_16; // @[IDU.scala 340:16]
  assign dpi_rf_17 = Registers_io_regs_17; // @[IDU.scala 341:16]
  assign dpi_rf_18 = Registers_io_regs_18; // @[IDU.scala 342:16]
  assign dpi_rf_19 = Registers_io_regs_19; // @[IDU.scala 343:16]
  assign dpi_rf_20 = Registers_io_regs_20; // @[IDU.scala 344:16]
  assign dpi_rf_21 = Registers_io_regs_21; // @[IDU.scala 345:16]
  assign dpi_rf_22 = Registers_io_regs_22; // @[IDU.scala 346:16]
  assign dpi_rf_23 = Registers_io_regs_23; // @[IDU.scala 347:16]
  assign dpi_rf_24 = Registers_io_regs_24; // @[IDU.scala 348:16]
  assign dpi_rf_25 = Registers_io_regs_25; // @[IDU.scala 349:16]
  assign dpi_rf_26 = Registers_io_regs_26; // @[IDU.scala 350:16]
  assign dpi_rf_27 = Registers_io_regs_27; // @[IDU.scala 351:16]
  assign dpi_rf_28 = Registers_io_regs_28; // @[IDU.scala 352:16]
  assign dpi_rf_29 = Registers_io_regs_29; // @[IDU.scala 353:16]
  assign dpi_rf_30 = Registers_io_regs_30; // @[IDU.scala 354:16]
  assign dpi_rf_31 = Registers_io_regs_31; // @[IDU.scala 355:16]
  assign dpi_csr_0 = CSR_io_csrs_0; // @[IDU.scala 358:16]
  assign dpi_csr_1 = CSR_io_csrs_1; // @[IDU.scala 359:16]
  assign dpi_csr_2 = CSR_io_csrs_2; // @[IDU.scala 360:16]
  assign dpi_csr_3 = CSR_io_csrs_3; // @[IDU.scala 361:16]
  assign dpi_csr_4 = CSR_io_csrs_4; // @[IDU.scala 362:16]
  assign dpi_inst = io_rf_bus_wb_inst; // @[IDU.scala 356:16]
  assign dpi_pc = {{32'd0}, io_rf_bus_wb_pc}; // @[IDU.scala 357:16]
  assign dpi_eval = {{31'd0}, eval}; // @[IDU.scala 363:16]
  always @(posedge clock) begin
    if (reset) begin // @[IDU.scala 31:28]
      ds_valid <= 1'h0; // @[IDU.scala 31:28]
    end else if (br_taken_cancel & io_ds_allowin) begin // @[IDU.scala 58:42]
      ds_valid <= 1'h0; // @[IDU.scala 59:14]
    end else if (io_ds_allowin) begin // @[IDU.scala 60:29]
      ds_valid <= io_fs_to_ds_valid; // @[IDU.scala 61:14]
    end
    if (reset) begin // @[IDU.scala 33:28]
      fd_bus_r_inst <= 32'h0; // @[IDU.scala 33:28]
    end else if (io_fs_to_ds_valid & io_ds_allowin) begin // @[IDU.scala 64:44]
      fd_bus_r_inst <= io_fd_bus_inst; // @[IDU.scala 65:14]
    end
    if (reset) begin // @[IDU.scala 33:28]
      fd_bus_r_pc <= 32'h0; // @[IDU.scala 33:28]
    end else if (io_fs_to_ds_valid & io_ds_allowin) begin // @[IDU.scala 64:44]
      fd_bus_r_pc <= io_fd_bus_pc; // @[IDU.scala 65:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ds_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  fd_bus_r_inst = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  fd_bus_r_pc = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RS(
  input   io_sel_negative,
  input   io_sel_positive,
  input   io_sel_double_negative,
  input   io_sel_double_positive,
  input   io_x,
  input   io_x_sub,
  output  io_p
);
  wire  _io_p_T_2 = ~(io_sel_negative & ~io_x); // @[RS.scala 17:11]
  wire  _io_p_T_6 = _io_p_T_2 & ~(io_sel_double_negative & ~io_x_sub); // @[RS.scala 18:9]
  wire  _io_p_T_9 = _io_p_T_6 & ~(io_sel_positive & io_x); // @[RS.scala 19:9]
  wire  _io_p_T_12 = _io_p_T_9 & ~(io_sel_double_positive & io_x_sub); // @[RS.scala 20:9]
  assign io_p = ~_io_p_T_12; // @[RS.scala 17:9]
endmodule
module BOOTH_S(
  output       io_sel_negative,
  output       io_sel_positive,
  output       io_sel_double_negative,
  output       io_sel_double_positive,
  output       io_cout,
  input  [2:0] io_src
);
  wire  y_add = io_src[2]; // @[BOOTH_S.scala 15:23]
  wire  y = io_src[1]; // @[BOOTH_S.scala 16:23]
  wire  y_sub = io_src[0]; // @[BOOTH_S.scala 17:23]
  wire  _io_sel_negative_T = ~y_sub; // @[BOOTH_S.scala 18:37]
  wire  _io_sel_negative_T_2 = ~y; // @[BOOTH_S.scala 18:46]
  wire  _io_sel_negative_T_4 = y & ~y_sub | ~y & y_sub; // @[BOOTH_S.scala 18:44]
  wire  _io_sel_negative_T_5 = y_add & (y & ~y_sub | ~y & y_sub); // @[BOOTH_S.scala 18:30]
  wire  _io_sel_positive_T = ~y_add; // @[BOOTH_S.scala 19:24]
  wire  _io_sel_double_negative_T_3 = y_add & _io_sel_negative_T_2 & _io_sel_negative_T; // @[BOOTH_S.scala 20:42]
  assign io_sel_negative = y_add & (y & ~y_sub | ~y & y_sub); // @[BOOTH_S.scala 18:30]
  assign io_sel_positive = ~y_add & _io_sel_negative_T_4; // @[BOOTH_S.scala 19:31]
  assign io_sel_double_negative = y_add & _io_sel_negative_T_2 & _io_sel_negative_T; // @[BOOTH_S.scala 20:42]
  assign io_sel_double_positive = _io_sel_positive_T & y & y_sub; // @[BOOTH_S.scala 21:42]
  assign io_cout = _io_sel_double_negative_T_3 | _io_sel_negative_T_5; // @[BOOTH_S.scala 22:38]
endmodule
module BOOTH_gen(
  input  [131:0] io_x,
  input  [2:0]   io_y,
  output [131:0] io_out,
  output         io_cout
);
  wire  RS_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_1_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_1_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_1_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_1_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_1_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_1_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_1_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_2_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_2_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_2_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_2_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_2_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_2_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_2_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_3_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_3_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_3_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_3_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_3_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_3_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_3_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_4_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_4_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_4_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_4_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_4_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_4_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_4_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_5_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_5_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_5_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_5_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_5_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_5_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_5_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_6_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_6_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_6_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_6_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_6_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_6_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_6_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_7_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_7_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_7_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_7_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_7_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_7_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_7_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_8_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_8_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_8_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_8_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_8_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_8_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_8_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_9_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_9_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_9_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_9_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_9_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_9_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_9_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_10_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_10_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_10_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_10_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_10_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_10_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_10_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_11_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_11_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_11_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_11_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_11_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_11_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_11_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_12_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_12_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_12_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_12_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_12_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_12_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_12_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_13_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_13_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_13_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_13_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_13_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_13_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_13_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_14_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_14_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_14_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_14_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_14_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_14_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_14_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_15_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_15_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_15_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_15_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_15_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_15_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_15_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_16_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_16_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_16_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_16_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_16_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_16_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_16_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_17_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_17_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_17_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_17_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_17_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_17_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_17_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_18_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_18_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_18_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_18_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_18_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_18_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_18_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_19_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_19_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_19_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_19_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_19_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_19_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_19_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_20_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_20_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_20_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_20_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_20_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_20_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_20_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_21_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_21_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_21_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_21_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_21_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_21_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_21_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_22_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_22_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_22_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_22_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_22_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_22_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_22_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_23_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_23_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_23_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_23_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_23_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_23_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_23_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_24_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_24_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_24_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_24_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_24_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_24_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_24_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_25_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_25_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_25_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_25_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_25_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_25_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_25_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_26_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_26_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_26_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_26_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_26_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_26_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_26_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_27_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_27_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_27_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_27_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_27_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_27_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_27_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_28_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_28_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_28_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_28_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_28_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_28_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_28_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_29_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_29_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_29_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_29_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_29_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_29_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_29_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_30_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_30_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_30_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_30_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_30_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_30_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_30_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_31_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_31_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_31_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_31_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_31_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_31_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_31_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_32_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_32_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_32_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_32_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_32_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_32_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_32_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_33_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_33_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_33_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_33_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_33_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_33_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_33_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_34_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_34_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_34_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_34_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_34_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_34_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_34_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_35_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_35_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_35_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_35_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_35_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_35_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_35_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_36_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_36_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_36_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_36_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_36_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_36_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_36_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_37_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_37_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_37_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_37_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_37_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_37_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_37_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_38_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_38_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_38_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_38_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_38_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_38_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_38_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_39_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_39_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_39_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_39_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_39_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_39_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_39_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_40_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_40_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_40_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_40_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_40_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_40_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_40_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_41_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_41_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_41_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_41_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_41_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_41_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_41_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_42_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_42_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_42_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_42_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_42_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_42_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_42_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_43_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_43_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_43_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_43_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_43_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_43_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_43_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_44_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_44_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_44_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_44_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_44_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_44_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_44_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_45_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_45_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_45_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_45_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_45_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_45_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_45_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_46_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_46_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_46_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_46_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_46_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_46_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_46_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_47_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_47_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_47_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_47_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_47_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_47_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_47_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_48_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_48_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_48_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_48_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_48_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_48_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_48_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_49_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_49_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_49_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_49_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_49_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_49_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_49_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_50_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_50_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_50_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_50_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_50_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_50_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_50_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_51_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_51_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_51_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_51_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_51_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_51_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_51_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_52_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_52_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_52_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_52_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_52_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_52_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_52_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_53_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_53_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_53_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_53_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_53_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_53_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_53_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_54_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_54_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_54_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_54_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_54_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_54_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_54_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_55_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_55_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_55_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_55_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_55_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_55_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_55_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_56_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_56_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_56_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_56_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_56_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_56_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_56_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_57_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_57_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_57_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_57_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_57_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_57_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_57_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_58_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_58_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_58_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_58_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_58_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_58_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_58_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_59_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_59_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_59_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_59_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_59_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_59_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_59_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_60_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_60_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_60_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_60_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_60_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_60_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_60_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_61_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_61_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_61_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_61_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_61_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_61_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_61_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_62_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_62_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_62_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_62_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_62_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_62_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_62_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_63_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_63_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_63_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_63_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_63_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_63_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_63_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_64_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_64_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_64_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_64_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_64_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_64_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_64_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_65_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_65_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_65_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_65_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_65_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_65_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_65_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_66_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_66_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_66_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_66_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_66_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_66_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_66_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_67_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_67_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_67_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_67_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_67_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_67_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_67_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_68_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_68_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_68_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_68_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_68_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_68_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_68_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_69_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_69_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_69_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_69_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_69_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_69_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_69_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_70_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_70_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_70_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_70_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_70_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_70_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_70_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_71_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_71_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_71_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_71_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_71_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_71_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_71_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_72_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_72_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_72_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_72_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_72_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_72_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_72_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_73_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_73_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_73_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_73_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_73_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_73_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_73_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_74_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_74_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_74_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_74_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_74_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_74_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_74_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_75_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_75_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_75_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_75_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_75_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_75_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_75_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_76_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_76_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_76_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_76_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_76_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_76_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_76_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_77_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_77_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_77_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_77_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_77_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_77_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_77_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_78_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_78_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_78_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_78_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_78_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_78_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_78_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_79_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_79_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_79_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_79_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_79_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_79_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_79_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_80_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_80_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_80_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_80_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_80_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_80_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_80_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_81_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_81_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_81_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_81_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_81_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_81_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_81_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_82_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_82_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_82_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_82_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_82_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_82_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_82_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_83_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_83_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_83_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_83_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_83_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_83_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_83_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_84_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_84_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_84_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_84_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_84_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_84_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_84_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_85_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_85_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_85_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_85_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_85_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_85_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_85_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_86_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_86_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_86_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_86_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_86_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_86_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_86_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_87_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_87_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_87_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_87_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_87_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_87_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_87_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_88_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_88_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_88_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_88_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_88_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_88_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_88_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_89_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_89_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_89_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_89_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_89_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_89_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_89_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_90_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_90_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_90_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_90_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_90_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_90_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_90_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_91_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_91_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_91_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_91_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_91_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_91_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_91_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_92_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_92_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_92_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_92_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_92_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_92_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_92_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_93_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_93_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_93_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_93_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_93_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_93_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_93_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_94_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_94_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_94_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_94_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_94_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_94_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_94_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_95_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_95_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_95_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_95_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_95_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_95_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_95_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_96_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_96_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_96_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_96_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_96_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_96_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_96_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_97_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_97_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_97_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_97_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_97_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_97_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_97_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_98_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_98_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_98_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_98_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_98_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_98_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_98_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_99_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_99_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_99_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_99_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_99_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_99_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_99_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_100_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_100_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_100_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_100_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_100_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_100_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_100_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_101_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_101_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_101_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_101_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_101_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_101_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_101_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_102_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_102_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_102_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_102_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_102_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_102_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_102_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_103_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_103_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_103_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_103_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_103_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_103_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_103_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_104_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_104_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_104_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_104_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_104_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_104_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_104_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_105_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_105_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_105_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_105_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_105_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_105_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_105_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_106_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_106_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_106_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_106_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_106_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_106_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_106_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_107_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_107_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_107_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_107_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_107_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_107_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_107_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_108_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_108_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_108_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_108_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_108_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_108_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_108_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_109_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_109_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_109_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_109_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_109_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_109_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_109_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_110_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_110_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_110_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_110_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_110_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_110_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_110_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_111_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_111_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_111_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_111_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_111_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_111_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_111_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_112_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_112_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_112_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_112_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_112_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_112_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_112_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_113_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_113_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_113_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_113_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_113_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_113_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_113_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_114_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_114_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_114_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_114_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_114_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_114_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_114_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_115_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_115_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_115_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_115_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_115_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_115_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_115_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_116_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_116_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_116_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_116_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_116_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_116_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_116_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_117_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_117_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_117_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_117_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_117_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_117_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_117_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_118_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_118_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_118_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_118_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_118_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_118_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_118_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_119_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_119_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_119_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_119_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_119_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_119_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_119_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_120_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_120_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_120_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_120_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_120_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_120_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_120_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_121_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_121_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_121_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_121_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_121_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_121_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_121_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_122_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_122_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_122_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_122_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_122_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_122_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_122_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_123_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_123_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_123_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_123_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_123_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_123_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_123_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_124_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_124_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_124_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_124_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_124_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_124_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_124_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_125_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_125_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_125_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_125_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_125_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_125_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_125_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_126_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_126_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_126_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_126_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_126_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_126_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_126_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_127_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_127_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_127_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_127_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_127_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_127_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_127_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_128_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_128_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_128_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_128_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_128_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_128_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_128_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_129_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_129_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_129_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_129_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_129_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_129_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_129_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_130_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_130_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_130_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_130_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_130_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_130_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_130_io_p; // @[BOOTH_gen.scala 16:42]
  wire  RS_131_io_sel_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_131_io_sel_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_131_io_sel_double_negative; // @[BOOTH_gen.scala 16:42]
  wire  RS_131_io_sel_double_positive; // @[BOOTH_gen.scala 16:42]
  wire  RS_131_io_x; // @[BOOTH_gen.scala 16:42]
  wire  RS_131_io_x_sub; // @[BOOTH_gen.scala 16:42]
  wire  RS_131_io_p; // @[BOOTH_gen.scala 16:42]
  wire  BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 17:21]
  wire  BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 17:21]
  wire  BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 17:21]
  wire  BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 17:21]
  wire  BOOTH_S_io_cout; // @[BOOTH_gen.scala 17:21]
  wire [2:0] BOOTH_S_io_src; // @[BOOTH_gen.scala 17:21]
  wire  r_1_p = RS_1_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_0_p = RS_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_3_p = RS_3_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_2_p = RS_2_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_5_p = RS_5_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_4_p = RS_4_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_7_p = RS_7_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_6_p = RS_6_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [7:0] io_out_lo_lo_lo_lo = {r_7_p,r_6_p,r_5_p,r_4_p,r_3_p,r_2_p,r_1_p,r_0_p}; // @[Cat.scala 31:58]
  wire  r_9_p = RS_9_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_8_p = RS_8_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_11_p = RS_11_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_10_p = RS_10_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_13_p = RS_13_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_12_p = RS_12_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_15_p = RS_15_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_14_p = RS_14_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_17_p = RS_17_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_16_p = RS_16_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_19_p = RS_19_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_18_p = RS_18_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_21_p = RS_21_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_20_p = RS_20_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_23_p = RS_23_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_22_p = RS_22_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [7:0] io_out_lo_lo_hi_lo = {r_23_p,r_22_p,r_21_p,r_20_p,r_19_p,r_18_p,r_17_p,r_16_p}; // @[Cat.scala 31:58]
  wire  r_25_p = RS_25_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_24_p = RS_24_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_27_p = RS_27_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_26_p = RS_26_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_29_p = RS_29_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_28_p = RS_28_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_32_p = RS_32_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_31_p = RS_31_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_30_p = RS_30_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [16:0] io_out_lo_lo_hi = {r_32_p,r_31_p,r_30_p,r_29_p,r_28_p,r_27_p,r_26_p,r_25_p,r_24_p,io_out_lo_lo_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] io_out_lo_lo = {io_out_lo_lo_hi,r_15_p,r_14_p,r_13_p,r_12_p,r_11_p,r_10_p,r_9_p,r_8_p,io_out_lo_lo_lo_lo}; // @[Cat.scala 31:58]
  wire  r_34_p = RS_34_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_33_p = RS_33_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_36_p = RS_36_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_35_p = RS_35_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_38_p = RS_38_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_37_p = RS_37_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_40_p = RS_40_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_39_p = RS_39_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [7:0] io_out_lo_hi_lo_lo = {r_40_p,r_39_p,r_38_p,r_37_p,r_36_p,r_35_p,r_34_p,r_33_p}; // @[Cat.scala 31:58]
  wire  r_42_p = RS_42_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_41_p = RS_41_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_44_p = RS_44_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_43_p = RS_43_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_46_p = RS_46_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_45_p = RS_45_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_48_p = RS_48_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_47_p = RS_47_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_50_p = RS_50_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_49_p = RS_49_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_52_p = RS_52_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_51_p = RS_51_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_54_p = RS_54_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_53_p = RS_53_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_56_p = RS_56_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_55_p = RS_55_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [7:0] io_out_lo_hi_hi_lo = {r_56_p,r_55_p,r_54_p,r_53_p,r_52_p,r_51_p,r_50_p,r_49_p}; // @[Cat.scala 31:58]
  wire  r_58_p = RS_58_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_57_p = RS_57_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_60_p = RS_60_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_59_p = RS_59_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_62_p = RS_62_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_61_p = RS_61_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_65_p = RS_65_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_64_p = RS_64_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_63_p = RS_63_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [16:0] io_out_lo_hi_hi = {r_65_p,r_64_p,r_63_p,r_62_p,r_61_p,r_60_p,r_59_p,r_58_p,r_57_p,io_out_lo_hi_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] io_out_lo_hi = {io_out_lo_hi_hi,r_48_p,r_47_p,r_46_p,r_45_p,r_44_p,r_43_p,r_42_p,r_41_p,io_out_lo_hi_lo_lo
    }; // @[Cat.scala 31:58]
  wire [65:0] io_out_lo = {io_out_lo_hi,io_out_lo_lo}; // @[Cat.scala 31:58]
  wire  r_67_p = RS_67_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_66_p = RS_66_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_69_p = RS_69_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_68_p = RS_68_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_71_p = RS_71_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_70_p = RS_70_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_73_p = RS_73_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_72_p = RS_72_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [7:0] io_out_hi_lo_lo_lo = {r_73_p,r_72_p,r_71_p,r_70_p,r_69_p,r_68_p,r_67_p,r_66_p}; // @[Cat.scala 31:58]
  wire  r_75_p = RS_75_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_74_p = RS_74_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_77_p = RS_77_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_76_p = RS_76_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_79_p = RS_79_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_78_p = RS_78_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_81_p = RS_81_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_80_p = RS_80_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_83_p = RS_83_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_82_p = RS_82_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_85_p = RS_85_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_84_p = RS_84_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_87_p = RS_87_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_86_p = RS_86_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_89_p = RS_89_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_88_p = RS_88_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [7:0] io_out_hi_lo_hi_lo = {r_89_p,r_88_p,r_87_p,r_86_p,r_85_p,r_84_p,r_83_p,r_82_p}; // @[Cat.scala 31:58]
  wire  r_91_p = RS_91_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_90_p = RS_90_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_93_p = RS_93_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_92_p = RS_92_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_95_p = RS_95_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_94_p = RS_94_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_98_p = RS_98_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_97_p = RS_97_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_96_p = RS_96_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [16:0] io_out_hi_lo_hi = {r_98_p,r_97_p,r_96_p,r_95_p,r_94_p,r_93_p,r_92_p,r_91_p,r_90_p,io_out_hi_lo_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] io_out_hi_lo = {io_out_hi_lo_hi,r_81_p,r_80_p,r_79_p,r_78_p,r_77_p,r_76_p,r_75_p,r_74_p,io_out_hi_lo_lo_lo
    }; // @[Cat.scala 31:58]
  wire  r_100_p = RS_100_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_99_p = RS_99_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_102_p = RS_102_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_101_p = RS_101_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_104_p = RS_104_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_103_p = RS_103_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_106_p = RS_106_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_105_p = RS_105_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [7:0] io_out_hi_hi_lo_lo = {r_106_p,r_105_p,r_104_p,r_103_p,r_102_p,r_101_p,r_100_p,r_99_p}; // @[Cat.scala 31:58]
  wire  r_108_p = RS_108_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_107_p = RS_107_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_110_p = RS_110_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_109_p = RS_109_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_112_p = RS_112_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_111_p = RS_111_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_114_p = RS_114_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_113_p = RS_113_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_116_p = RS_116_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_115_p = RS_115_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_118_p = RS_118_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_117_p = RS_117_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_120_p = RS_120_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_119_p = RS_119_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_122_p = RS_122_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_121_p = RS_121_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [7:0] io_out_hi_hi_hi_lo = {r_122_p,r_121_p,r_120_p,r_119_p,r_118_p,r_117_p,r_116_p,r_115_p}; // @[Cat.scala 31:58]
  wire  r_124_p = RS_124_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_123_p = RS_123_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_126_p = RS_126_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_125_p = RS_125_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_128_p = RS_128_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_127_p = RS_127_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_131_p = RS_131_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_130_p = RS_130_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire  r_129_p = RS_129_io_p; // @[BOOTH_gen.scala 16:{20,20}]
  wire [16:0] io_out_hi_hi_hi = {r_131_p,r_130_p,r_129_p,r_128_p,r_127_p,r_126_p,r_125_p,r_124_p,r_123_p,
    io_out_hi_hi_hi_lo}; // @[Cat.scala 31:58]
  wire [32:0] io_out_hi_hi = {io_out_hi_hi_hi,r_114_p,r_113_p,r_112_p,r_111_p,r_110_p,r_109_p,r_108_p,r_107_p,
    io_out_hi_hi_lo_lo}; // @[Cat.scala 31:58]
  wire [65:0] io_out_hi = {io_out_hi_hi,io_out_hi_lo}; // @[Cat.scala 31:58]
  RS RS ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_io_sel_negative),
    .io_sel_positive(RS_io_sel_positive),
    .io_sel_double_negative(RS_io_sel_double_negative),
    .io_sel_double_positive(RS_io_sel_double_positive),
    .io_x(RS_io_x),
    .io_x_sub(RS_io_x_sub),
    .io_p(RS_io_p)
  );
  RS RS_1 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_1_io_sel_negative),
    .io_sel_positive(RS_1_io_sel_positive),
    .io_sel_double_negative(RS_1_io_sel_double_negative),
    .io_sel_double_positive(RS_1_io_sel_double_positive),
    .io_x(RS_1_io_x),
    .io_x_sub(RS_1_io_x_sub),
    .io_p(RS_1_io_p)
  );
  RS RS_2 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_2_io_sel_negative),
    .io_sel_positive(RS_2_io_sel_positive),
    .io_sel_double_negative(RS_2_io_sel_double_negative),
    .io_sel_double_positive(RS_2_io_sel_double_positive),
    .io_x(RS_2_io_x),
    .io_x_sub(RS_2_io_x_sub),
    .io_p(RS_2_io_p)
  );
  RS RS_3 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_3_io_sel_negative),
    .io_sel_positive(RS_3_io_sel_positive),
    .io_sel_double_negative(RS_3_io_sel_double_negative),
    .io_sel_double_positive(RS_3_io_sel_double_positive),
    .io_x(RS_3_io_x),
    .io_x_sub(RS_3_io_x_sub),
    .io_p(RS_3_io_p)
  );
  RS RS_4 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_4_io_sel_negative),
    .io_sel_positive(RS_4_io_sel_positive),
    .io_sel_double_negative(RS_4_io_sel_double_negative),
    .io_sel_double_positive(RS_4_io_sel_double_positive),
    .io_x(RS_4_io_x),
    .io_x_sub(RS_4_io_x_sub),
    .io_p(RS_4_io_p)
  );
  RS RS_5 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_5_io_sel_negative),
    .io_sel_positive(RS_5_io_sel_positive),
    .io_sel_double_negative(RS_5_io_sel_double_negative),
    .io_sel_double_positive(RS_5_io_sel_double_positive),
    .io_x(RS_5_io_x),
    .io_x_sub(RS_5_io_x_sub),
    .io_p(RS_5_io_p)
  );
  RS RS_6 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_6_io_sel_negative),
    .io_sel_positive(RS_6_io_sel_positive),
    .io_sel_double_negative(RS_6_io_sel_double_negative),
    .io_sel_double_positive(RS_6_io_sel_double_positive),
    .io_x(RS_6_io_x),
    .io_x_sub(RS_6_io_x_sub),
    .io_p(RS_6_io_p)
  );
  RS RS_7 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_7_io_sel_negative),
    .io_sel_positive(RS_7_io_sel_positive),
    .io_sel_double_negative(RS_7_io_sel_double_negative),
    .io_sel_double_positive(RS_7_io_sel_double_positive),
    .io_x(RS_7_io_x),
    .io_x_sub(RS_7_io_x_sub),
    .io_p(RS_7_io_p)
  );
  RS RS_8 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_8_io_sel_negative),
    .io_sel_positive(RS_8_io_sel_positive),
    .io_sel_double_negative(RS_8_io_sel_double_negative),
    .io_sel_double_positive(RS_8_io_sel_double_positive),
    .io_x(RS_8_io_x),
    .io_x_sub(RS_8_io_x_sub),
    .io_p(RS_8_io_p)
  );
  RS RS_9 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_9_io_sel_negative),
    .io_sel_positive(RS_9_io_sel_positive),
    .io_sel_double_negative(RS_9_io_sel_double_negative),
    .io_sel_double_positive(RS_9_io_sel_double_positive),
    .io_x(RS_9_io_x),
    .io_x_sub(RS_9_io_x_sub),
    .io_p(RS_9_io_p)
  );
  RS RS_10 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_10_io_sel_negative),
    .io_sel_positive(RS_10_io_sel_positive),
    .io_sel_double_negative(RS_10_io_sel_double_negative),
    .io_sel_double_positive(RS_10_io_sel_double_positive),
    .io_x(RS_10_io_x),
    .io_x_sub(RS_10_io_x_sub),
    .io_p(RS_10_io_p)
  );
  RS RS_11 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_11_io_sel_negative),
    .io_sel_positive(RS_11_io_sel_positive),
    .io_sel_double_negative(RS_11_io_sel_double_negative),
    .io_sel_double_positive(RS_11_io_sel_double_positive),
    .io_x(RS_11_io_x),
    .io_x_sub(RS_11_io_x_sub),
    .io_p(RS_11_io_p)
  );
  RS RS_12 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_12_io_sel_negative),
    .io_sel_positive(RS_12_io_sel_positive),
    .io_sel_double_negative(RS_12_io_sel_double_negative),
    .io_sel_double_positive(RS_12_io_sel_double_positive),
    .io_x(RS_12_io_x),
    .io_x_sub(RS_12_io_x_sub),
    .io_p(RS_12_io_p)
  );
  RS RS_13 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_13_io_sel_negative),
    .io_sel_positive(RS_13_io_sel_positive),
    .io_sel_double_negative(RS_13_io_sel_double_negative),
    .io_sel_double_positive(RS_13_io_sel_double_positive),
    .io_x(RS_13_io_x),
    .io_x_sub(RS_13_io_x_sub),
    .io_p(RS_13_io_p)
  );
  RS RS_14 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_14_io_sel_negative),
    .io_sel_positive(RS_14_io_sel_positive),
    .io_sel_double_negative(RS_14_io_sel_double_negative),
    .io_sel_double_positive(RS_14_io_sel_double_positive),
    .io_x(RS_14_io_x),
    .io_x_sub(RS_14_io_x_sub),
    .io_p(RS_14_io_p)
  );
  RS RS_15 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_15_io_sel_negative),
    .io_sel_positive(RS_15_io_sel_positive),
    .io_sel_double_negative(RS_15_io_sel_double_negative),
    .io_sel_double_positive(RS_15_io_sel_double_positive),
    .io_x(RS_15_io_x),
    .io_x_sub(RS_15_io_x_sub),
    .io_p(RS_15_io_p)
  );
  RS RS_16 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_16_io_sel_negative),
    .io_sel_positive(RS_16_io_sel_positive),
    .io_sel_double_negative(RS_16_io_sel_double_negative),
    .io_sel_double_positive(RS_16_io_sel_double_positive),
    .io_x(RS_16_io_x),
    .io_x_sub(RS_16_io_x_sub),
    .io_p(RS_16_io_p)
  );
  RS RS_17 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_17_io_sel_negative),
    .io_sel_positive(RS_17_io_sel_positive),
    .io_sel_double_negative(RS_17_io_sel_double_negative),
    .io_sel_double_positive(RS_17_io_sel_double_positive),
    .io_x(RS_17_io_x),
    .io_x_sub(RS_17_io_x_sub),
    .io_p(RS_17_io_p)
  );
  RS RS_18 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_18_io_sel_negative),
    .io_sel_positive(RS_18_io_sel_positive),
    .io_sel_double_negative(RS_18_io_sel_double_negative),
    .io_sel_double_positive(RS_18_io_sel_double_positive),
    .io_x(RS_18_io_x),
    .io_x_sub(RS_18_io_x_sub),
    .io_p(RS_18_io_p)
  );
  RS RS_19 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_19_io_sel_negative),
    .io_sel_positive(RS_19_io_sel_positive),
    .io_sel_double_negative(RS_19_io_sel_double_negative),
    .io_sel_double_positive(RS_19_io_sel_double_positive),
    .io_x(RS_19_io_x),
    .io_x_sub(RS_19_io_x_sub),
    .io_p(RS_19_io_p)
  );
  RS RS_20 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_20_io_sel_negative),
    .io_sel_positive(RS_20_io_sel_positive),
    .io_sel_double_negative(RS_20_io_sel_double_negative),
    .io_sel_double_positive(RS_20_io_sel_double_positive),
    .io_x(RS_20_io_x),
    .io_x_sub(RS_20_io_x_sub),
    .io_p(RS_20_io_p)
  );
  RS RS_21 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_21_io_sel_negative),
    .io_sel_positive(RS_21_io_sel_positive),
    .io_sel_double_negative(RS_21_io_sel_double_negative),
    .io_sel_double_positive(RS_21_io_sel_double_positive),
    .io_x(RS_21_io_x),
    .io_x_sub(RS_21_io_x_sub),
    .io_p(RS_21_io_p)
  );
  RS RS_22 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_22_io_sel_negative),
    .io_sel_positive(RS_22_io_sel_positive),
    .io_sel_double_negative(RS_22_io_sel_double_negative),
    .io_sel_double_positive(RS_22_io_sel_double_positive),
    .io_x(RS_22_io_x),
    .io_x_sub(RS_22_io_x_sub),
    .io_p(RS_22_io_p)
  );
  RS RS_23 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_23_io_sel_negative),
    .io_sel_positive(RS_23_io_sel_positive),
    .io_sel_double_negative(RS_23_io_sel_double_negative),
    .io_sel_double_positive(RS_23_io_sel_double_positive),
    .io_x(RS_23_io_x),
    .io_x_sub(RS_23_io_x_sub),
    .io_p(RS_23_io_p)
  );
  RS RS_24 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_24_io_sel_negative),
    .io_sel_positive(RS_24_io_sel_positive),
    .io_sel_double_negative(RS_24_io_sel_double_negative),
    .io_sel_double_positive(RS_24_io_sel_double_positive),
    .io_x(RS_24_io_x),
    .io_x_sub(RS_24_io_x_sub),
    .io_p(RS_24_io_p)
  );
  RS RS_25 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_25_io_sel_negative),
    .io_sel_positive(RS_25_io_sel_positive),
    .io_sel_double_negative(RS_25_io_sel_double_negative),
    .io_sel_double_positive(RS_25_io_sel_double_positive),
    .io_x(RS_25_io_x),
    .io_x_sub(RS_25_io_x_sub),
    .io_p(RS_25_io_p)
  );
  RS RS_26 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_26_io_sel_negative),
    .io_sel_positive(RS_26_io_sel_positive),
    .io_sel_double_negative(RS_26_io_sel_double_negative),
    .io_sel_double_positive(RS_26_io_sel_double_positive),
    .io_x(RS_26_io_x),
    .io_x_sub(RS_26_io_x_sub),
    .io_p(RS_26_io_p)
  );
  RS RS_27 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_27_io_sel_negative),
    .io_sel_positive(RS_27_io_sel_positive),
    .io_sel_double_negative(RS_27_io_sel_double_negative),
    .io_sel_double_positive(RS_27_io_sel_double_positive),
    .io_x(RS_27_io_x),
    .io_x_sub(RS_27_io_x_sub),
    .io_p(RS_27_io_p)
  );
  RS RS_28 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_28_io_sel_negative),
    .io_sel_positive(RS_28_io_sel_positive),
    .io_sel_double_negative(RS_28_io_sel_double_negative),
    .io_sel_double_positive(RS_28_io_sel_double_positive),
    .io_x(RS_28_io_x),
    .io_x_sub(RS_28_io_x_sub),
    .io_p(RS_28_io_p)
  );
  RS RS_29 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_29_io_sel_negative),
    .io_sel_positive(RS_29_io_sel_positive),
    .io_sel_double_negative(RS_29_io_sel_double_negative),
    .io_sel_double_positive(RS_29_io_sel_double_positive),
    .io_x(RS_29_io_x),
    .io_x_sub(RS_29_io_x_sub),
    .io_p(RS_29_io_p)
  );
  RS RS_30 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_30_io_sel_negative),
    .io_sel_positive(RS_30_io_sel_positive),
    .io_sel_double_negative(RS_30_io_sel_double_negative),
    .io_sel_double_positive(RS_30_io_sel_double_positive),
    .io_x(RS_30_io_x),
    .io_x_sub(RS_30_io_x_sub),
    .io_p(RS_30_io_p)
  );
  RS RS_31 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_31_io_sel_negative),
    .io_sel_positive(RS_31_io_sel_positive),
    .io_sel_double_negative(RS_31_io_sel_double_negative),
    .io_sel_double_positive(RS_31_io_sel_double_positive),
    .io_x(RS_31_io_x),
    .io_x_sub(RS_31_io_x_sub),
    .io_p(RS_31_io_p)
  );
  RS RS_32 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_32_io_sel_negative),
    .io_sel_positive(RS_32_io_sel_positive),
    .io_sel_double_negative(RS_32_io_sel_double_negative),
    .io_sel_double_positive(RS_32_io_sel_double_positive),
    .io_x(RS_32_io_x),
    .io_x_sub(RS_32_io_x_sub),
    .io_p(RS_32_io_p)
  );
  RS RS_33 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_33_io_sel_negative),
    .io_sel_positive(RS_33_io_sel_positive),
    .io_sel_double_negative(RS_33_io_sel_double_negative),
    .io_sel_double_positive(RS_33_io_sel_double_positive),
    .io_x(RS_33_io_x),
    .io_x_sub(RS_33_io_x_sub),
    .io_p(RS_33_io_p)
  );
  RS RS_34 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_34_io_sel_negative),
    .io_sel_positive(RS_34_io_sel_positive),
    .io_sel_double_negative(RS_34_io_sel_double_negative),
    .io_sel_double_positive(RS_34_io_sel_double_positive),
    .io_x(RS_34_io_x),
    .io_x_sub(RS_34_io_x_sub),
    .io_p(RS_34_io_p)
  );
  RS RS_35 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_35_io_sel_negative),
    .io_sel_positive(RS_35_io_sel_positive),
    .io_sel_double_negative(RS_35_io_sel_double_negative),
    .io_sel_double_positive(RS_35_io_sel_double_positive),
    .io_x(RS_35_io_x),
    .io_x_sub(RS_35_io_x_sub),
    .io_p(RS_35_io_p)
  );
  RS RS_36 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_36_io_sel_negative),
    .io_sel_positive(RS_36_io_sel_positive),
    .io_sel_double_negative(RS_36_io_sel_double_negative),
    .io_sel_double_positive(RS_36_io_sel_double_positive),
    .io_x(RS_36_io_x),
    .io_x_sub(RS_36_io_x_sub),
    .io_p(RS_36_io_p)
  );
  RS RS_37 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_37_io_sel_negative),
    .io_sel_positive(RS_37_io_sel_positive),
    .io_sel_double_negative(RS_37_io_sel_double_negative),
    .io_sel_double_positive(RS_37_io_sel_double_positive),
    .io_x(RS_37_io_x),
    .io_x_sub(RS_37_io_x_sub),
    .io_p(RS_37_io_p)
  );
  RS RS_38 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_38_io_sel_negative),
    .io_sel_positive(RS_38_io_sel_positive),
    .io_sel_double_negative(RS_38_io_sel_double_negative),
    .io_sel_double_positive(RS_38_io_sel_double_positive),
    .io_x(RS_38_io_x),
    .io_x_sub(RS_38_io_x_sub),
    .io_p(RS_38_io_p)
  );
  RS RS_39 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_39_io_sel_negative),
    .io_sel_positive(RS_39_io_sel_positive),
    .io_sel_double_negative(RS_39_io_sel_double_negative),
    .io_sel_double_positive(RS_39_io_sel_double_positive),
    .io_x(RS_39_io_x),
    .io_x_sub(RS_39_io_x_sub),
    .io_p(RS_39_io_p)
  );
  RS RS_40 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_40_io_sel_negative),
    .io_sel_positive(RS_40_io_sel_positive),
    .io_sel_double_negative(RS_40_io_sel_double_negative),
    .io_sel_double_positive(RS_40_io_sel_double_positive),
    .io_x(RS_40_io_x),
    .io_x_sub(RS_40_io_x_sub),
    .io_p(RS_40_io_p)
  );
  RS RS_41 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_41_io_sel_negative),
    .io_sel_positive(RS_41_io_sel_positive),
    .io_sel_double_negative(RS_41_io_sel_double_negative),
    .io_sel_double_positive(RS_41_io_sel_double_positive),
    .io_x(RS_41_io_x),
    .io_x_sub(RS_41_io_x_sub),
    .io_p(RS_41_io_p)
  );
  RS RS_42 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_42_io_sel_negative),
    .io_sel_positive(RS_42_io_sel_positive),
    .io_sel_double_negative(RS_42_io_sel_double_negative),
    .io_sel_double_positive(RS_42_io_sel_double_positive),
    .io_x(RS_42_io_x),
    .io_x_sub(RS_42_io_x_sub),
    .io_p(RS_42_io_p)
  );
  RS RS_43 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_43_io_sel_negative),
    .io_sel_positive(RS_43_io_sel_positive),
    .io_sel_double_negative(RS_43_io_sel_double_negative),
    .io_sel_double_positive(RS_43_io_sel_double_positive),
    .io_x(RS_43_io_x),
    .io_x_sub(RS_43_io_x_sub),
    .io_p(RS_43_io_p)
  );
  RS RS_44 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_44_io_sel_negative),
    .io_sel_positive(RS_44_io_sel_positive),
    .io_sel_double_negative(RS_44_io_sel_double_negative),
    .io_sel_double_positive(RS_44_io_sel_double_positive),
    .io_x(RS_44_io_x),
    .io_x_sub(RS_44_io_x_sub),
    .io_p(RS_44_io_p)
  );
  RS RS_45 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_45_io_sel_negative),
    .io_sel_positive(RS_45_io_sel_positive),
    .io_sel_double_negative(RS_45_io_sel_double_negative),
    .io_sel_double_positive(RS_45_io_sel_double_positive),
    .io_x(RS_45_io_x),
    .io_x_sub(RS_45_io_x_sub),
    .io_p(RS_45_io_p)
  );
  RS RS_46 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_46_io_sel_negative),
    .io_sel_positive(RS_46_io_sel_positive),
    .io_sel_double_negative(RS_46_io_sel_double_negative),
    .io_sel_double_positive(RS_46_io_sel_double_positive),
    .io_x(RS_46_io_x),
    .io_x_sub(RS_46_io_x_sub),
    .io_p(RS_46_io_p)
  );
  RS RS_47 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_47_io_sel_negative),
    .io_sel_positive(RS_47_io_sel_positive),
    .io_sel_double_negative(RS_47_io_sel_double_negative),
    .io_sel_double_positive(RS_47_io_sel_double_positive),
    .io_x(RS_47_io_x),
    .io_x_sub(RS_47_io_x_sub),
    .io_p(RS_47_io_p)
  );
  RS RS_48 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_48_io_sel_negative),
    .io_sel_positive(RS_48_io_sel_positive),
    .io_sel_double_negative(RS_48_io_sel_double_negative),
    .io_sel_double_positive(RS_48_io_sel_double_positive),
    .io_x(RS_48_io_x),
    .io_x_sub(RS_48_io_x_sub),
    .io_p(RS_48_io_p)
  );
  RS RS_49 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_49_io_sel_negative),
    .io_sel_positive(RS_49_io_sel_positive),
    .io_sel_double_negative(RS_49_io_sel_double_negative),
    .io_sel_double_positive(RS_49_io_sel_double_positive),
    .io_x(RS_49_io_x),
    .io_x_sub(RS_49_io_x_sub),
    .io_p(RS_49_io_p)
  );
  RS RS_50 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_50_io_sel_negative),
    .io_sel_positive(RS_50_io_sel_positive),
    .io_sel_double_negative(RS_50_io_sel_double_negative),
    .io_sel_double_positive(RS_50_io_sel_double_positive),
    .io_x(RS_50_io_x),
    .io_x_sub(RS_50_io_x_sub),
    .io_p(RS_50_io_p)
  );
  RS RS_51 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_51_io_sel_negative),
    .io_sel_positive(RS_51_io_sel_positive),
    .io_sel_double_negative(RS_51_io_sel_double_negative),
    .io_sel_double_positive(RS_51_io_sel_double_positive),
    .io_x(RS_51_io_x),
    .io_x_sub(RS_51_io_x_sub),
    .io_p(RS_51_io_p)
  );
  RS RS_52 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_52_io_sel_negative),
    .io_sel_positive(RS_52_io_sel_positive),
    .io_sel_double_negative(RS_52_io_sel_double_negative),
    .io_sel_double_positive(RS_52_io_sel_double_positive),
    .io_x(RS_52_io_x),
    .io_x_sub(RS_52_io_x_sub),
    .io_p(RS_52_io_p)
  );
  RS RS_53 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_53_io_sel_negative),
    .io_sel_positive(RS_53_io_sel_positive),
    .io_sel_double_negative(RS_53_io_sel_double_negative),
    .io_sel_double_positive(RS_53_io_sel_double_positive),
    .io_x(RS_53_io_x),
    .io_x_sub(RS_53_io_x_sub),
    .io_p(RS_53_io_p)
  );
  RS RS_54 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_54_io_sel_negative),
    .io_sel_positive(RS_54_io_sel_positive),
    .io_sel_double_negative(RS_54_io_sel_double_negative),
    .io_sel_double_positive(RS_54_io_sel_double_positive),
    .io_x(RS_54_io_x),
    .io_x_sub(RS_54_io_x_sub),
    .io_p(RS_54_io_p)
  );
  RS RS_55 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_55_io_sel_negative),
    .io_sel_positive(RS_55_io_sel_positive),
    .io_sel_double_negative(RS_55_io_sel_double_negative),
    .io_sel_double_positive(RS_55_io_sel_double_positive),
    .io_x(RS_55_io_x),
    .io_x_sub(RS_55_io_x_sub),
    .io_p(RS_55_io_p)
  );
  RS RS_56 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_56_io_sel_negative),
    .io_sel_positive(RS_56_io_sel_positive),
    .io_sel_double_negative(RS_56_io_sel_double_negative),
    .io_sel_double_positive(RS_56_io_sel_double_positive),
    .io_x(RS_56_io_x),
    .io_x_sub(RS_56_io_x_sub),
    .io_p(RS_56_io_p)
  );
  RS RS_57 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_57_io_sel_negative),
    .io_sel_positive(RS_57_io_sel_positive),
    .io_sel_double_negative(RS_57_io_sel_double_negative),
    .io_sel_double_positive(RS_57_io_sel_double_positive),
    .io_x(RS_57_io_x),
    .io_x_sub(RS_57_io_x_sub),
    .io_p(RS_57_io_p)
  );
  RS RS_58 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_58_io_sel_negative),
    .io_sel_positive(RS_58_io_sel_positive),
    .io_sel_double_negative(RS_58_io_sel_double_negative),
    .io_sel_double_positive(RS_58_io_sel_double_positive),
    .io_x(RS_58_io_x),
    .io_x_sub(RS_58_io_x_sub),
    .io_p(RS_58_io_p)
  );
  RS RS_59 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_59_io_sel_negative),
    .io_sel_positive(RS_59_io_sel_positive),
    .io_sel_double_negative(RS_59_io_sel_double_negative),
    .io_sel_double_positive(RS_59_io_sel_double_positive),
    .io_x(RS_59_io_x),
    .io_x_sub(RS_59_io_x_sub),
    .io_p(RS_59_io_p)
  );
  RS RS_60 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_60_io_sel_negative),
    .io_sel_positive(RS_60_io_sel_positive),
    .io_sel_double_negative(RS_60_io_sel_double_negative),
    .io_sel_double_positive(RS_60_io_sel_double_positive),
    .io_x(RS_60_io_x),
    .io_x_sub(RS_60_io_x_sub),
    .io_p(RS_60_io_p)
  );
  RS RS_61 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_61_io_sel_negative),
    .io_sel_positive(RS_61_io_sel_positive),
    .io_sel_double_negative(RS_61_io_sel_double_negative),
    .io_sel_double_positive(RS_61_io_sel_double_positive),
    .io_x(RS_61_io_x),
    .io_x_sub(RS_61_io_x_sub),
    .io_p(RS_61_io_p)
  );
  RS RS_62 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_62_io_sel_negative),
    .io_sel_positive(RS_62_io_sel_positive),
    .io_sel_double_negative(RS_62_io_sel_double_negative),
    .io_sel_double_positive(RS_62_io_sel_double_positive),
    .io_x(RS_62_io_x),
    .io_x_sub(RS_62_io_x_sub),
    .io_p(RS_62_io_p)
  );
  RS RS_63 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_63_io_sel_negative),
    .io_sel_positive(RS_63_io_sel_positive),
    .io_sel_double_negative(RS_63_io_sel_double_negative),
    .io_sel_double_positive(RS_63_io_sel_double_positive),
    .io_x(RS_63_io_x),
    .io_x_sub(RS_63_io_x_sub),
    .io_p(RS_63_io_p)
  );
  RS RS_64 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_64_io_sel_negative),
    .io_sel_positive(RS_64_io_sel_positive),
    .io_sel_double_negative(RS_64_io_sel_double_negative),
    .io_sel_double_positive(RS_64_io_sel_double_positive),
    .io_x(RS_64_io_x),
    .io_x_sub(RS_64_io_x_sub),
    .io_p(RS_64_io_p)
  );
  RS RS_65 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_65_io_sel_negative),
    .io_sel_positive(RS_65_io_sel_positive),
    .io_sel_double_negative(RS_65_io_sel_double_negative),
    .io_sel_double_positive(RS_65_io_sel_double_positive),
    .io_x(RS_65_io_x),
    .io_x_sub(RS_65_io_x_sub),
    .io_p(RS_65_io_p)
  );
  RS RS_66 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_66_io_sel_negative),
    .io_sel_positive(RS_66_io_sel_positive),
    .io_sel_double_negative(RS_66_io_sel_double_negative),
    .io_sel_double_positive(RS_66_io_sel_double_positive),
    .io_x(RS_66_io_x),
    .io_x_sub(RS_66_io_x_sub),
    .io_p(RS_66_io_p)
  );
  RS RS_67 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_67_io_sel_negative),
    .io_sel_positive(RS_67_io_sel_positive),
    .io_sel_double_negative(RS_67_io_sel_double_negative),
    .io_sel_double_positive(RS_67_io_sel_double_positive),
    .io_x(RS_67_io_x),
    .io_x_sub(RS_67_io_x_sub),
    .io_p(RS_67_io_p)
  );
  RS RS_68 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_68_io_sel_negative),
    .io_sel_positive(RS_68_io_sel_positive),
    .io_sel_double_negative(RS_68_io_sel_double_negative),
    .io_sel_double_positive(RS_68_io_sel_double_positive),
    .io_x(RS_68_io_x),
    .io_x_sub(RS_68_io_x_sub),
    .io_p(RS_68_io_p)
  );
  RS RS_69 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_69_io_sel_negative),
    .io_sel_positive(RS_69_io_sel_positive),
    .io_sel_double_negative(RS_69_io_sel_double_negative),
    .io_sel_double_positive(RS_69_io_sel_double_positive),
    .io_x(RS_69_io_x),
    .io_x_sub(RS_69_io_x_sub),
    .io_p(RS_69_io_p)
  );
  RS RS_70 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_70_io_sel_negative),
    .io_sel_positive(RS_70_io_sel_positive),
    .io_sel_double_negative(RS_70_io_sel_double_negative),
    .io_sel_double_positive(RS_70_io_sel_double_positive),
    .io_x(RS_70_io_x),
    .io_x_sub(RS_70_io_x_sub),
    .io_p(RS_70_io_p)
  );
  RS RS_71 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_71_io_sel_negative),
    .io_sel_positive(RS_71_io_sel_positive),
    .io_sel_double_negative(RS_71_io_sel_double_negative),
    .io_sel_double_positive(RS_71_io_sel_double_positive),
    .io_x(RS_71_io_x),
    .io_x_sub(RS_71_io_x_sub),
    .io_p(RS_71_io_p)
  );
  RS RS_72 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_72_io_sel_negative),
    .io_sel_positive(RS_72_io_sel_positive),
    .io_sel_double_negative(RS_72_io_sel_double_negative),
    .io_sel_double_positive(RS_72_io_sel_double_positive),
    .io_x(RS_72_io_x),
    .io_x_sub(RS_72_io_x_sub),
    .io_p(RS_72_io_p)
  );
  RS RS_73 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_73_io_sel_negative),
    .io_sel_positive(RS_73_io_sel_positive),
    .io_sel_double_negative(RS_73_io_sel_double_negative),
    .io_sel_double_positive(RS_73_io_sel_double_positive),
    .io_x(RS_73_io_x),
    .io_x_sub(RS_73_io_x_sub),
    .io_p(RS_73_io_p)
  );
  RS RS_74 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_74_io_sel_negative),
    .io_sel_positive(RS_74_io_sel_positive),
    .io_sel_double_negative(RS_74_io_sel_double_negative),
    .io_sel_double_positive(RS_74_io_sel_double_positive),
    .io_x(RS_74_io_x),
    .io_x_sub(RS_74_io_x_sub),
    .io_p(RS_74_io_p)
  );
  RS RS_75 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_75_io_sel_negative),
    .io_sel_positive(RS_75_io_sel_positive),
    .io_sel_double_negative(RS_75_io_sel_double_negative),
    .io_sel_double_positive(RS_75_io_sel_double_positive),
    .io_x(RS_75_io_x),
    .io_x_sub(RS_75_io_x_sub),
    .io_p(RS_75_io_p)
  );
  RS RS_76 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_76_io_sel_negative),
    .io_sel_positive(RS_76_io_sel_positive),
    .io_sel_double_negative(RS_76_io_sel_double_negative),
    .io_sel_double_positive(RS_76_io_sel_double_positive),
    .io_x(RS_76_io_x),
    .io_x_sub(RS_76_io_x_sub),
    .io_p(RS_76_io_p)
  );
  RS RS_77 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_77_io_sel_negative),
    .io_sel_positive(RS_77_io_sel_positive),
    .io_sel_double_negative(RS_77_io_sel_double_negative),
    .io_sel_double_positive(RS_77_io_sel_double_positive),
    .io_x(RS_77_io_x),
    .io_x_sub(RS_77_io_x_sub),
    .io_p(RS_77_io_p)
  );
  RS RS_78 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_78_io_sel_negative),
    .io_sel_positive(RS_78_io_sel_positive),
    .io_sel_double_negative(RS_78_io_sel_double_negative),
    .io_sel_double_positive(RS_78_io_sel_double_positive),
    .io_x(RS_78_io_x),
    .io_x_sub(RS_78_io_x_sub),
    .io_p(RS_78_io_p)
  );
  RS RS_79 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_79_io_sel_negative),
    .io_sel_positive(RS_79_io_sel_positive),
    .io_sel_double_negative(RS_79_io_sel_double_negative),
    .io_sel_double_positive(RS_79_io_sel_double_positive),
    .io_x(RS_79_io_x),
    .io_x_sub(RS_79_io_x_sub),
    .io_p(RS_79_io_p)
  );
  RS RS_80 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_80_io_sel_negative),
    .io_sel_positive(RS_80_io_sel_positive),
    .io_sel_double_negative(RS_80_io_sel_double_negative),
    .io_sel_double_positive(RS_80_io_sel_double_positive),
    .io_x(RS_80_io_x),
    .io_x_sub(RS_80_io_x_sub),
    .io_p(RS_80_io_p)
  );
  RS RS_81 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_81_io_sel_negative),
    .io_sel_positive(RS_81_io_sel_positive),
    .io_sel_double_negative(RS_81_io_sel_double_negative),
    .io_sel_double_positive(RS_81_io_sel_double_positive),
    .io_x(RS_81_io_x),
    .io_x_sub(RS_81_io_x_sub),
    .io_p(RS_81_io_p)
  );
  RS RS_82 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_82_io_sel_negative),
    .io_sel_positive(RS_82_io_sel_positive),
    .io_sel_double_negative(RS_82_io_sel_double_negative),
    .io_sel_double_positive(RS_82_io_sel_double_positive),
    .io_x(RS_82_io_x),
    .io_x_sub(RS_82_io_x_sub),
    .io_p(RS_82_io_p)
  );
  RS RS_83 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_83_io_sel_negative),
    .io_sel_positive(RS_83_io_sel_positive),
    .io_sel_double_negative(RS_83_io_sel_double_negative),
    .io_sel_double_positive(RS_83_io_sel_double_positive),
    .io_x(RS_83_io_x),
    .io_x_sub(RS_83_io_x_sub),
    .io_p(RS_83_io_p)
  );
  RS RS_84 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_84_io_sel_negative),
    .io_sel_positive(RS_84_io_sel_positive),
    .io_sel_double_negative(RS_84_io_sel_double_negative),
    .io_sel_double_positive(RS_84_io_sel_double_positive),
    .io_x(RS_84_io_x),
    .io_x_sub(RS_84_io_x_sub),
    .io_p(RS_84_io_p)
  );
  RS RS_85 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_85_io_sel_negative),
    .io_sel_positive(RS_85_io_sel_positive),
    .io_sel_double_negative(RS_85_io_sel_double_negative),
    .io_sel_double_positive(RS_85_io_sel_double_positive),
    .io_x(RS_85_io_x),
    .io_x_sub(RS_85_io_x_sub),
    .io_p(RS_85_io_p)
  );
  RS RS_86 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_86_io_sel_negative),
    .io_sel_positive(RS_86_io_sel_positive),
    .io_sel_double_negative(RS_86_io_sel_double_negative),
    .io_sel_double_positive(RS_86_io_sel_double_positive),
    .io_x(RS_86_io_x),
    .io_x_sub(RS_86_io_x_sub),
    .io_p(RS_86_io_p)
  );
  RS RS_87 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_87_io_sel_negative),
    .io_sel_positive(RS_87_io_sel_positive),
    .io_sel_double_negative(RS_87_io_sel_double_negative),
    .io_sel_double_positive(RS_87_io_sel_double_positive),
    .io_x(RS_87_io_x),
    .io_x_sub(RS_87_io_x_sub),
    .io_p(RS_87_io_p)
  );
  RS RS_88 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_88_io_sel_negative),
    .io_sel_positive(RS_88_io_sel_positive),
    .io_sel_double_negative(RS_88_io_sel_double_negative),
    .io_sel_double_positive(RS_88_io_sel_double_positive),
    .io_x(RS_88_io_x),
    .io_x_sub(RS_88_io_x_sub),
    .io_p(RS_88_io_p)
  );
  RS RS_89 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_89_io_sel_negative),
    .io_sel_positive(RS_89_io_sel_positive),
    .io_sel_double_negative(RS_89_io_sel_double_negative),
    .io_sel_double_positive(RS_89_io_sel_double_positive),
    .io_x(RS_89_io_x),
    .io_x_sub(RS_89_io_x_sub),
    .io_p(RS_89_io_p)
  );
  RS RS_90 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_90_io_sel_negative),
    .io_sel_positive(RS_90_io_sel_positive),
    .io_sel_double_negative(RS_90_io_sel_double_negative),
    .io_sel_double_positive(RS_90_io_sel_double_positive),
    .io_x(RS_90_io_x),
    .io_x_sub(RS_90_io_x_sub),
    .io_p(RS_90_io_p)
  );
  RS RS_91 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_91_io_sel_negative),
    .io_sel_positive(RS_91_io_sel_positive),
    .io_sel_double_negative(RS_91_io_sel_double_negative),
    .io_sel_double_positive(RS_91_io_sel_double_positive),
    .io_x(RS_91_io_x),
    .io_x_sub(RS_91_io_x_sub),
    .io_p(RS_91_io_p)
  );
  RS RS_92 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_92_io_sel_negative),
    .io_sel_positive(RS_92_io_sel_positive),
    .io_sel_double_negative(RS_92_io_sel_double_negative),
    .io_sel_double_positive(RS_92_io_sel_double_positive),
    .io_x(RS_92_io_x),
    .io_x_sub(RS_92_io_x_sub),
    .io_p(RS_92_io_p)
  );
  RS RS_93 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_93_io_sel_negative),
    .io_sel_positive(RS_93_io_sel_positive),
    .io_sel_double_negative(RS_93_io_sel_double_negative),
    .io_sel_double_positive(RS_93_io_sel_double_positive),
    .io_x(RS_93_io_x),
    .io_x_sub(RS_93_io_x_sub),
    .io_p(RS_93_io_p)
  );
  RS RS_94 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_94_io_sel_negative),
    .io_sel_positive(RS_94_io_sel_positive),
    .io_sel_double_negative(RS_94_io_sel_double_negative),
    .io_sel_double_positive(RS_94_io_sel_double_positive),
    .io_x(RS_94_io_x),
    .io_x_sub(RS_94_io_x_sub),
    .io_p(RS_94_io_p)
  );
  RS RS_95 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_95_io_sel_negative),
    .io_sel_positive(RS_95_io_sel_positive),
    .io_sel_double_negative(RS_95_io_sel_double_negative),
    .io_sel_double_positive(RS_95_io_sel_double_positive),
    .io_x(RS_95_io_x),
    .io_x_sub(RS_95_io_x_sub),
    .io_p(RS_95_io_p)
  );
  RS RS_96 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_96_io_sel_negative),
    .io_sel_positive(RS_96_io_sel_positive),
    .io_sel_double_negative(RS_96_io_sel_double_negative),
    .io_sel_double_positive(RS_96_io_sel_double_positive),
    .io_x(RS_96_io_x),
    .io_x_sub(RS_96_io_x_sub),
    .io_p(RS_96_io_p)
  );
  RS RS_97 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_97_io_sel_negative),
    .io_sel_positive(RS_97_io_sel_positive),
    .io_sel_double_negative(RS_97_io_sel_double_negative),
    .io_sel_double_positive(RS_97_io_sel_double_positive),
    .io_x(RS_97_io_x),
    .io_x_sub(RS_97_io_x_sub),
    .io_p(RS_97_io_p)
  );
  RS RS_98 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_98_io_sel_negative),
    .io_sel_positive(RS_98_io_sel_positive),
    .io_sel_double_negative(RS_98_io_sel_double_negative),
    .io_sel_double_positive(RS_98_io_sel_double_positive),
    .io_x(RS_98_io_x),
    .io_x_sub(RS_98_io_x_sub),
    .io_p(RS_98_io_p)
  );
  RS RS_99 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_99_io_sel_negative),
    .io_sel_positive(RS_99_io_sel_positive),
    .io_sel_double_negative(RS_99_io_sel_double_negative),
    .io_sel_double_positive(RS_99_io_sel_double_positive),
    .io_x(RS_99_io_x),
    .io_x_sub(RS_99_io_x_sub),
    .io_p(RS_99_io_p)
  );
  RS RS_100 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_100_io_sel_negative),
    .io_sel_positive(RS_100_io_sel_positive),
    .io_sel_double_negative(RS_100_io_sel_double_negative),
    .io_sel_double_positive(RS_100_io_sel_double_positive),
    .io_x(RS_100_io_x),
    .io_x_sub(RS_100_io_x_sub),
    .io_p(RS_100_io_p)
  );
  RS RS_101 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_101_io_sel_negative),
    .io_sel_positive(RS_101_io_sel_positive),
    .io_sel_double_negative(RS_101_io_sel_double_negative),
    .io_sel_double_positive(RS_101_io_sel_double_positive),
    .io_x(RS_101_io_x),
    .io_x_sub(RS_101_io_x_sub),
    .io_p(RS_101_io_p)
  );
  RS RS_102 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_102_io_sel_negative),
    .io_sel_positive(RS_102_io_sel_positive),
    .io_sel_double_negative(RS_102_io_sel_double_negative),
    .io_sel_double_positive(RS_102_io_sel_double_positive),
    .io_x(RS_102_io_x),
    .io_x_sub(RS_102_io_x_sub),
    .io_p(RS_102_io_p)
  );
  RS RS_103 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_103_io_sel_negative),
    .io_sel_positive(RS_103_io_sel_positive),
    .io_sel_double_negative(RS_103_io_sel_double_negative),
    .io_sel_double_positive(RS_103_io_sel_double_positive),
    .io_x(RS_103_io_x),
    .io_x_sub(RS_103_io_x_sub),
    .io_p(RS_103_io_p)
  );
  RS RS_104 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_104_io_sel_negative),
    .io_sel_positive(RS_104_io_sel_positive),
    .io_sel_double_negative(RS_104_io_sel_double_negative),
    .io_sel_double_positive(RS_104_io_sel_double_positive),
    .io_x(RS_104_io_x),
    .io_x_sub(RS_104_io_x_sub),
    .io_p(RS_104_io_p)
  );
  RS RS_105 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_105_io_sel_negative),
    .io_sel_positive(RS_105_io_sel_positive),
    .io_sel_double_negative(RS_105_io_sel_double_negative),
    .io_sel_double_positive(RS_105_io_sel_double_positive),
    .io_x(RS_105_io_x),
    .io_x_sub(RS_105_io_x_sub),
    .io_p(RS_105_io_p)
  );
  RS RS_106 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_106_io_sel_negative),
    .io_sel_positive(RS_106_io_sel_positive),
    .io_sel_double_negative(RS_106_io_sel_double_negative),
    .io_sel_double_positive(RS_106_io_sel_double_positive),
    .io_x(RS_106_io_x),
    .io_x_sub(RS_106_io_x_sub),
    .io_p(RS_106_io_p)
  );
  RS RS_107 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_107_io_sel_negative),
    .io_sel_positive(RS_107_io_sel_positive),
    .io_sel_double_negative(RS_107_io_sel_double_negative),
    .io_sel_double_positive(RS_107_io_sel_double_positive),
    .io_x(RS_107_io_x),
    .io_x_sub(RS_107_io_x_sub),
    .io_p(RS_107_io_p)
  );
  RS RS_108 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_108_io_sel_negative),
    .io_sel_positive(RS_108_io_sel_positive),
    .io_sel_double_negative(RS_108_io_sel_double_negative),
    .io_sel_double_positive(RS_108_io_sel_double_positive),
    .io_x(RS_108_io_x),
    .io_x_sub(RS_108_io_x_sub),
    .io_p(RS_108_io_p)
  );
  RS RS_109 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_109_io_sel_negative),
    .io_sel_positive(RS_109_io_sel_positive),
    .io_sel_double_negative(RS_109_io_sel_double_negative),
    .io_sel_double_positive(RS_109_io_sel_double_positive),
    .io_x(RS_109_io_x),
    .io_x_sub(RS_109_io_x_sub),
    .io_p(RS_109_io_p)
  );
  RS RS_110 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_110_io_sel_negative),
    .io_sel_positive(RS_110_io_sel_positive),
    .io_sel_double_negative(RS_110_io_sel_double_negative),
    .io_sel_double_positive(RS_110_io_sel_double_positive),
    .io_x(RS_110_io_x),
    .io_x_sub(RS_110_io_x_sub),
    .io_p(RS_110_io_p)
  );
  RS RS_111 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_111_io_sel_negative),
    .io_sel_positive(RS_111_io_sel_positive),
    .io_sel_double_negative(RS_111_io_sel_double_negative),
    .io_sel_double_positive(RS_111_io_sel_double_positive),
    .io_x(RS_111_io_x),
    .io_x_sub(RS_111_io_x_sub),
    .io_p(RS_111_io_p)
  );
  RS RS_112 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_112_io_sel_negative),
    .io_sel_positive(RS_112_io_sel_positive),
    .io_sel_double_negative(RS_112_io_sel_double_negative),
    .io_sel_double_positive(RS_112_io_sel_double_positive),
    .io_x(RS_112_io_x),
    .io_x_sub(RS_112_io_x_sub),
    .io_p(RS_112_io_p)
  );
  RS RS_113 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_113_io_sel_negative),
    .io_sel_positive(RS_113_io_sel_positive),
    .io_sel_double_negative(RS_113_io_sel_double_negative),
    .io_sel_double_positive(RS_113_io_sel_double_positive),
    .io_x(RS_113_io_x),
    .io_x_sub(RS_113_io_x_sub),
    .io_p(RS_113_io_p)
  );
  RS RS_114 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_114_io_sel_negative),
    .io_sel_positive(RS_114_io_sel_positive),
    .io_sel_double_negative(RS_114_io_sel_double_negative),
    .io_sel_double_positive(RS_114_io_sel_double_positive),
    .io_x(RS_114_io_x),
    .io_x_sub(RS_114_io_x_sub),
    .io_p(RS_114_io_p)
  );
  RS RS_115 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_115_io_sel_negative),
    .io_sel_positive(RS_115_io_sel_positive),
    .io_sel_double_negative(RS_115_io_sel_double_negative),
    .io_sel_double_positive(RS_115_io_sel_double_positive),
    .io_x(RS_115_io_x),
    .io_x_sub(RS_115_io_x_sub),
    .io_p(RS_115_io_p)
  );
  RS RS_116 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_116_io_sel_negative),
    .io_sel_positive(RS_116_io_sel_positive),
    .io_sel_double_negative(RS_116_io_sel_double_negative),
    .io_sel_double_positive(RS_116_io_sel_double_positive),
    .io_x(RS_116_io_x),
    .io_x_sub(RS_116_io_x_sub),
    .io_p(RS_116_io_p)
  );
  RS RS_117 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_117_io_sel_negative),
    .io_sel_positive(RS_117_io_sel_positive),
    .io_sel_double_negative(RS_117_io_sel_double_negative),
    .io_sel_double_positive(RS_117_io_sel_double_positive),
    .io_x(RS_117_io_x),
    .io_x_sub(RS_117_io_x_sub),
    .io_p(RS_117_io_p)
  );
  RS RS_118 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_118_io_sel_negative),
    .io_sel_positive(RS_118_io_sel_positive),
    .io_sel_double_negative(RS_118_io_sel_double_negative),
    .io_sel_double_positive(RS_118_io_sel_double_positive),
    .io_x(RS_118_io_x),
    .io_x_sub(RS_118_io_x_sub),
    .io_p(RS_118_io_p)
  );
  RS RS_119 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_119_io_sel_negative),
    .io_sel_positive(RS_119_io_sel_positive),
    .io_sel_double_negative(RS_119_io_sel_double_negative),
    .io_sel_double_positive(RS_119_io_sel_double_positive),
    .io_x(RS_119_io_x),
    .io_x_sub(RS_119_io_x_sub),
    .io_p(RS_119_io_p)
  );
  RS RS_120 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_120_io_sel_negative),
    .io_sel_positive(RS_120_io_sel_positive),
    .io_sel_double_negative(RS_120_io_sel_double_negative),
    .io_sel_double_positive(RS_120_io_sel_double_positive),
    .io_x(RS_120_io_x),
    .io_x_sub(RS_120_io_x_sub),
    .io_p(RS_120_io_p)
  );
  RS RS_121 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_121_io_sel_negative),
    .io_sel_positive(RS_121_io_sel_positive),
    .io_sel_double_negative(RS_121_io_sel_double_negative),
    .io_sel_double_positive(RS_121_io_sel_double_positive),
    .io_x(RS_121_io_x),
    .io_x_sub(RS_121_io_x_sub),
    .io_p(RS_121_io_p)
  );
  RS RS_122 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_122_io_sel_negative),
    .io_sel_positive(RS_122_io_sel_positive),
    .io_sel_double_negative(RS_122_io_sel_double_negative),
    .io_sel_double_positive(RS_122_io_sel_double_positive),
    .io_x(RS_122_io_x),
    .io_x_sub(RS_122_io_x_sub),
    .io_p(RS_122_io_p)
  );
  RS RS_123 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_123_io_sel_negative),
    .io_sel_positive(RS_123_io_sel_positive),
    .io_sel_double_negative(RS_123_io_sel_double_negative),
    .io_sel_double_positive(RS_123_io_sel_double_positive),
    .io_x(RS_123_io_x),
    .io_x_sub(RS_123_io_x_sub),
    .io_p(RS_123_io_p)
  );
  RS RS_124 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_124_io_sel_negative),
    .io_sel_positive(RS_124_io_sel_positive),
    .io_sel_double_negative(RS_124_io_sel_double_negative),
    .io_sel_double_positive(RS_124_io_sel_double_positive),
    .io_x(RS_124_io_x),
    .io_x_sub(RS_124_io_x_sub),
    .io_p(RS_124_io_p)
  );
  RS RS_125 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_125_io_sel_negative),
    .io_sel_positive(RS_125_io_sel_positive),
    .io_sel_double_negative(RS_125_io_sel_double_negative),
    .io_sel_double_positive(RS_125_io_sel_double_positive),
    .io_x(RS_125_io_x),
    .io_x_sub(RS_125_io_x_sub),
    .io_p(RS_125_io_p)
  );
  RS RS_126 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_126_io_sel_negative),
    .io_sel_positive(RS_126_io_sel_positive),
    .io_sel_double_negative(RS_126_io_sel_double_negative),
    .io_sel_double_positive(RS_126_io_sel_double_positive),
    .io_x(RS_126_io_x),
    .io_x_sub(RS_126_io_x_sub),
    .io_p(RS_126_io_p)
  );
  RS RS_127 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_127_io_sel_negative),
    .io_sel_positive(RS_127_io_sel_positive),
    .io_sel_double_negative(RS_127_io_sel_double_negative),
    .io_sel_double_positive(RS_127_io_sel_double_positive),
    .io_x(RS_127_io_x),
    .io_x_sub(RS_127_io_x_sub),
    .io_p(RS_127_io_p)
  );
  RS RS_128 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_128_io_sel_negative),
    .io_sel_positive(RS_128_io_sel_positive),
    .io_sel_double_negative(RS_128_io_sel_double_negative),
    .io_sel_double_positive(RS_128_io_sel_double_positive),
    .io_x(RS_128_io_x),
    .io_x_sub(RS_128_io_x_sub),
    .io_p(RS_128_io_p)
  );
  RS RS_129 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_129_io_sel_negative),
    .io_sel_positive(RS_129_io_sel_positive),
    .io_sel_double_negative(RS_129_io_sel_double_negative),
    .io_sel_double_positive(RS_129_io_sel_double_positive),
    .io_x(RS_129_io_x),
    .io_x_sub(RS_129_io_x_sub),
    .io_p(RS_129_io_p)
  );
  RS RS_130 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_130_io_sel_negative),
    .io_sel_positive(RS_130_io_sel_positive),
    .io_sel_double_negative(RS_130_io_sel_double_negative),
    .io_sel_double_positive(RS_130_io_sel_double_positive),
    .io_x(RS_130_io_x),
    .io_x_sub(RS_130_io_x_sub),
    .io_p(RS_130_io_p)
  );
  RS RS_131 ( // @[BOOTH_gen.scala 16:42]
    .io_sel_negative(RS_131_io_sel_negative),
    .io_sel_positive(RS_131_io_sel_positive),
    .io_sel_double_negative(RS_131_io_sel_double_negative),
    .io_sel_double_positive(RS_131_io_sel_double_positive),
    .io_x(RS_131_io_x),
    .io_x_sub(RS_131_io_x_sub),
    .io_p(RS_131_io_p)
  );
  BOOTH_S BOOTH_S ( // @[BOOTH_gen.scala 17:21]
    .io_sel_negative(BOOTH_S_io_sel_negative),
    .io_sel_positive(BOOTH_S_io_sel_positive),
    .io_sel_double_negative(BOOTH_S_io_sel_double_negative),
    .io_sel_double_positive(BOOTH_S_io_sel_double_positive),
    .io_cout(BOOTH_S_io_cout),
    .io_src(BOOTH_S_io_src)
  );
  assign io_out = {io_out_hi,io_out_lo}; // @[Cat.scala 31:58]
  assign io_cout = BOOTH_S_io_cout; // @[BOOTH_gen.scala 38:13]
  assign RS_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 23:23]
  assign RS_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 24:23]
  assign RS_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 25:30]
  assign RS_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 26:30]
  assign RS_io_x = io_x[0]; // @[BOOTH_gen.scala 21:16]
  assign RS_io_x_sub = 1'h0; // @[BOOTH_gen.scala 16:20 22:16]
  assign RS_1_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_1_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_1_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_1_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_1_io_x = io_x[1]; // @[BOOTH_gen.scala 29:20]
  assign RS_1_io_x_sub = io_x[0]; // @[BOOTH_gen.scala 30:24]
  assign RS_2_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_2_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_2_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_2_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_2_io_x = io_x[2]; // @[BOOTH_gen.scala 29:20]
  assign RS_2_io_x_sub = io_x[1]; // @[BOOTH_gen.scala 30:24]
  assign RS_3_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_3_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_3_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_3_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_3_io_x = io_x[3]; // @[BOOTH_gen.scala 29:20]
  assign RS_3_io_x_sub = io_x[2]; // @[BOOTH_gen.scala 30:24]
  assign RS_4_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_4_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_4_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_4_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_4_io_x = io_x[4]; // @[BOOTH_gen.scala 29:20]
  assign RS_4_io_x_sub = io_x[3]; // @[BOOTH_gen.scala 30:24]
  assign RS_5_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_5_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_5_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_5_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_5_io_x = io_x[5]; // @[BOOTH_gen.scala 29:20]
  assign RS_5_io_x_sub = io_x[4]; // @[BOOTH_gen.scala 30:24]
  assign RS_6_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_6_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_6_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_6_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_6_io_x = io_x[6]; // @[BOOTH_gen.scala 29:20]
  assign RS_6_io_x_sub = io_x[5]; // @[BOOTH_gen.scala 30:24]
  assign RS_7_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_7_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_7_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_7_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_7_io_x = io_x[7]; // @[BOOTH_gen.scala 29:20]
  assign RS_7_io_x_sub = io_x[6]; // @[BOOTH_gen.scala 30:24]
  assign RS_8_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_8_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_8_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_8_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_8_io_x = io_x[8]; // @[BOOTH_gen.scala 29:20]
  assign RS_8_io_x_sub = io_x[7]; // @[BOOTH_gen.scala 30:24]
  assign RS_9_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_9_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_9_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_9_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_9_io_x = io_x[9]; // @[BOOTH_gen.scala 29:20]
  assign RS_9_io_x_sub = io_x[8]; // @[BOOTH_gen.scala 30:24]
  assign RS_10_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_10_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_10_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_10_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_10_io_x = io_x[10]; // @[BOOTH_gen.scala 29:20]
  assign RS_10_io_x_sub = io_x[9]; // @[BOOTH_gen.scala 30:24]
  assign RS_11_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_11_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_11_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_11_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_11_io_x = io_x[11]; // @[BOOTH_gen.scala 29:20]
  assign RS_11_io_x_sub = io_x[10]; // @[BOOTH_gen.scala 30:24]
  assign RS_12_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_12_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_12_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_12_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_12_io_x = io_x[12]; // @[BOOTH_gen.scala 29:20]
  assign RS_12_io_x_sub = io_x[11]; // @[BOOTH_gen.scala 30:24]
  assign RS_13_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_13_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_13_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_13_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_13_io_x = io_x[13]; // @[BOOTH_gen.scala 29:20]
  assign RS_13_io_x_sub = io_x[12]; // @[BOOTH_gen.scala 30:24]
  assign RS_14_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_14_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_14_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_14_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_14_io_x = io_x[14]; // @[BOOTH_gen.scala 29:20]
  assign RS_14_io_x_sub = io_x[13]; // @[BOOTH_gen.scala 30:24]
  assign RS_15_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_15_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_15_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_15_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_15_io_x = io_x[15]; // @[BOOTH_gen.scala 29:20]
  assign RS_15_io_x_sub = io_x[14]; // @[BOOTH_gen.scala 30:24]
  assign RS_16_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_16_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_16_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_16_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_16_io_x = io_x[16]; // @[BOOTH_gen.scala 29:20]
  assign RS_16_io_x_sub = io_x[15]; // @[BOOTH_gen.scala 30:24]
  assign RS_17_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_17_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_17_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_17_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_17_io_x = io_x[17]; // @[BOOTH_gen.scala 29:20]
  assign RS_17_io_x_sub = io_x[16]; // @[BOOTH_gen.scala 30:24]
  assign RS_18_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_18_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_18_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_18_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_18_io_x = io_x[18]; // @[BOOTH_gen.scala 29:20]
  assign RS_18_io_x_sub = io_x[17]; // @[BOOTH_gen.scala 30:24]
  assign RS_19_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_19_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_19_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_19_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_19_io_x = io_x[19]; // @[BOOTH_gen.scala 29:20]
  assign RS_19_io_x_sub = io_x[18]; // @[BOOTH_gen.scala 30:24]
  assign RS_20_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_20_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_20_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_20_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_20_io_x = io_x[20]; // @[BOOTH_gen.scala 29:20]
  assign RS_20_io_x_sub = io_x[19]; // @[BOOTH_gen.scala 30:24]
  assign RS_21_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_21_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_21_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_21_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_21_io_x = io_x[21]; // @[BOOTH_gen.scala 29:20]
  assign RS_21_io_x_sub = io_x[20]; // @[BOOTH_gen.scala 30:24]
  assign RS_22_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_22_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_22_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_22_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_22_io_x = io_x[22]; // @[BOOTH_gen.scala 29:20]
  assign RS_22_io_x_sub = io_x[21]; // @[BOOTH_gen.scala 30:24]
  assign RS_23_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_23_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_23_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_23_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_23_io_x = io_x[23]; // @[BOOTH_gen.scala 29:20]
  assign RS_23_io_x_sub = io_x[22]; // @[BOOTH_gen.scala 30:24]
  assign RS_24_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_24_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_24_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_24_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_24_io_x = io_x[24]; // @[BOOTH_gen.scala 29:20]
  assign RS_24_io_x_sub = io_x[23]; // @[BOOTH_gen.scala 30:24]
  assign RS_25_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_25_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_25_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_25_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_25_io_x = io_x[25]; // @[BOOTH_gen.scala 29:20]
  assign RS_25_io_x_sub = io_x[24]; // @[BOOTH_gen.scala 30:24]
  assign RS_26_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_26_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_26_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_26_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_26_io_x = io_x[26]; // @[BOOTH_gen.scala 29:20]
  assign RS_26_io_x_sub = io_x[25]; // @[BOOTH_gen.scala 30:24]
  assign RS_27_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_27_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_27_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_27_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_27_io_x = io_x[27]; // @[BOOTH_gen.scala 29:20]
  assign RS_27_io_x_sub = io_x[26]; // @[BOOTH_gen.scala 30:24]
  assign RS_28_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_28_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_28_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_28_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_28_io_x = io_x[28]; // @[BOOTH_gen.scala 29:20]
  assign RS_28_io_x_sub = io_x[27]; // @[BOOTH_gen.scala 30:24]
  assign RS_29_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_29_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_29_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_29_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_29_io_x = io_x[29]; // @[BOOTH_gen.scala 29:20]
  assign RS_29_io_x_sub = io_x[28]; // @[BOOTH_gen.scala 30:24]
  assign RS_30_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_30_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_30_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_30_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_30_io_x = io_x[30]; // @[BOOTH_gen.scala 29:20]
  assign RS_30_io_x_sub = io_x[29]; // @[BOOTH_gen.scala 30:24]
  assign RS_31_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_31_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_31_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_31_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_31_io_x = io_x[31]; // @[BOOTH_gen.scala 29:20]
  assign RS_31_io_x_sub = io_x[30]; // @[BOOTH_gen.scala 30:24]
  assign RS_32_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_32_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_32_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_32_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_32_io_x = io_x[32]; // @[BOOTH_gen.scala 29:20]
  assign RS_32_io_x_sub = io_x[31]; // @[BOOTH_gen.scala 30:24]
  assign RS_33_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_33_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_33_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_33_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_33_io_x = io_x[33]; // @[BOOTH_gen.scala 29:20]
  assign RS_33_io_x_sub = io_x[32]; // @[BOOTH_gen.scala 30:24]
  assign RS_34_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_34_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_34_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_34_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_34_io_x = io_x[34]; // @[BOOTH_gen.scala 29:20]
  assign RS_34_io_x_sub = io_x[33]; // @[BOOTH_gen.scala 30:24]
  assign RS_35_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_35_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_35_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_35_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_35_io_x = io_x[35]; // @[BOOTH_gen.scala 29:20]
  assign RS_35_io_x_sub = io_x[34]; // @[BOOTH_gen.scala 30:24]
  assign RS_36_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_36_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_36_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_36_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_36_io_x = io_x[36]; // @[BOOTH_gen.scala 29:20]
  assign RS_36_io_x_sub = io_x[35]; // @[BOOTH_gen.scala 30:24]
  assign RS_37_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_37_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_37_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_37_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_37_io_x = io_x[37]; // @[BOOTH_gen.scala 29:20]
  assign RS_37_io_x_sub = io_x[36]; // @[BOOTH_gen.scala 30:24]
  assign RS_38_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_38_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_38_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_38_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_38_io_x = io_x[38]; // @[BOOTH_gen.scala 29:20]
  assign RS_38_io_x_sub = io_x[37]; // @[BOOTH_gen.scala 30:24]
  assign RS_39_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_39_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_39_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_39_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_39_io_x = io_x[39]; // @[BOOTH_gen.scala 29:20]
  assign RS_39_io_x_sub = io_x[38]; // @[BOOTH_gen.scala 30:24]
  assign RS_40_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_40_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_40_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_40_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_40_io_x = io_x[40]; // @[BOOTH_gen.scala 29:20]
  assign RS_40_io_x_sub = io_x[39]; // @[BOOTH_gen.scala 30:24]
  assign RS_41_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_41_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_41_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_41_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_41_io_x = io_x[41]; // @[BOOTH_gen.scala 29:20]
  assign RS_41_io_x_sub = io_x[40]; // @[BOOTH_gen.scala 30:24]
  assign RS_42_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_42_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_42_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_42_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_42_io_x = io_x[42]; // @[BOOTH_gen.scala 29:20]
  assign RS_42_io_x_sub = io_x[41]; // @[BOOTH_gen.scala 30:24]
  assign RS_43_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_43_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_43_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_43_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_43_io_x = io_x[43]; // @[BOOTH_gen.scala 29:20]
  assign RS_43_io_x_sub = io_x[42]; // @[BOOTH_gen.scala 30:24]
  assign RS_44_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_44_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_44_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_44_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_44_io_x = io_x[44]; // @[BOOTH_gen.scala 29:20]
  assign RS_44_io_x_sub = io_x[43]; // @[BOOTH_gen.scala 30:24]
  assign RS_45_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_45_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_45_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_45_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_45_io_x = io_x[45]; // @[BOOTH_gen.scala 29:20]
  assign RS_45_io_x_sub = io_x[44]; // @[BOOTH_gen.scala 30:24]
  assign RS_46_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_46_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_46_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_46_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_46_io_x = io_x[46]; // @[BOOTH_gen.scala 29:20]
  assign RS_46_io_x_sub = io_x[45]; // @[BOOTH_gen.scala 30:24]
  assign RS_47_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_47_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_47_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_47_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_47_io_x = io_x[47]; // @[BOOTH_gen.scala 29:20]
  assign RS_47_io_x_sub = io_x[46]; // @[BOOTH_gen.scala 30:24]
  assign RS_48_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_48_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_48_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_48_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_48_io_x = io_x[48]; // @[BOOTH_gen.scala 29:20]
  assign RS_48_io_x_sub = io_x[47]; // @[BOOTH_gen.scala 30:24]
  assign RS_49_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_49_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_49_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_49_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_49_io_x = io_x[49]; // @[BOOTH_gen.scala 29:20]
  assign RS_49_io_x_sub = io_x[48]; // @[BOOTH_gen.scala 30:24]
  assign RS_50_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_50_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_50_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_50_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_50_io_x = io_x[50]; // @[BOOTH_gen.scala 29:20]
  assign RS_50_io_x_sub = io_x[49]; // @[BOOTH_gen.scala 30:24]
  assign RS_51_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_51_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_51_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_51_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_51_io_x = io_x[51]; // @[BOOTH_gen.scala 29:20]
  assign RS_51_io_x_sub = io_x[50]; // @[BOOTH_gen.scala 30:24]
  assign RS_52_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_52_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_52_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_52_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_52_io_x = io_x[52]; // @[BOOTH_gen.scala 29:20]
  assign RS_52_io_x_sub = io_x[51]; // @[BOOTH_gen.scala 30:24]
  assign RS_53_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_53_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_53_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_53_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_53_io_x = io_x[53]; // @[BOOTH_gen.scala 29:20]
  assign RS_53_io_x_sub = io_x[52]; // @[BOOTH_gen.scala 30:24]
  assign RS_54_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_54_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_54_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_54_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_54_io_x = io_x[54]; // @[BOOTH_gen.scala 29:20]
  assign RS_54_io_x_sub = io_x[53]; // @[BOOTH_gen.scala 30:24]
  assign RS_55_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_55_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_55_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_55_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_55_io_x = io_x[55]; // @[BOOTH_gen.scala 29:20]
  assign RS_55_io_x_sub = io_x[54]; // @[BOOTH_gen.scala 30:24]
  assign RS_56_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_56_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_56_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_56_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_56_io_x = io_x[56]; // @[BOOTH_gen.scala 29:20]
  assign RS_56_io_x_sub = io_x[55]; // @[BOOTH_gen.scala 30:24]
  assign RS_57_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_57_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_57_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_57_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_57_io_x = io_x[57]; // @[BOOTH_gen.scala 29:20]
  assign RS_57_io_x_sub = io_x[56]; // @[BOOTH_gen.scala 30:24]
  assign RS_58_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_58_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_58_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_58_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_58_io_x = io_x[58]; // @[BOOTH_gen.scala 29:20]
  assign RS_58_io_x_sub = io_x[57]; // @[BOOTH_gen.scala 30:24]
  assign RS_59_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_59_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_59_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_59_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_59_io_x = io_x[59]; // @[BOOTH_gen.scala 29:20]
  assign RS_59_io_x_sub = io_x[58]; // @[BOOTH_gen.scala 30:24]
  assign RS_60_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_60_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_60_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_60_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_60_io_x = io_x[60]; // @[BOOTH_gen.scala 29:20]
  assign RS_60_io_x_sub = io_x[59]; // @[BOOTH_gen.scala 30:24]
  assign RS_61_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_61_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_61_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_61_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_61_io_x = io_x[61]; // @[BOOTH_gen.scala 29:20]
  assign RS_61_io_x_sub = io_x[60]; // @[BOOTH_gen.scala 30:24]
  assign RS_62_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_62_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_62_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_62_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_62_io_x = io_x[62]; // @[BOOTH_gen.scala 29:20]
  assign RS_62_io_x_sub = io_x[61]; // @[BOOTH_gen.scala 30:24]
  assign RS_63_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_63_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_63_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_63_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_63_io_x = io_x[63]; // @[BOOTH_gen.scala 29:20]
  assign RS_63_io_x_sub = io_x[62]; // @[BOOTH_gen.scala 30:24]
  assign RS_64_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_64_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_64_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_64_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_64_io_x = io_x[64]; // @[BOOTH_gen.scala 29:20]
  assign RS_64_io_x_sub = io_x[63]; // @[BOOTH_gen.scala 30:24]
  assign RS_65_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_65_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_65_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_65_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_65_io_x = io_x[65]; // @[BOOTH_gen.scala 29:20]
  assign RS_65_io_x_sub = io_x[64]; // @[BOOTH_gen.scala 30:24]
  assign RS_66_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_66_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_66_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_66_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_66_io_x = io_x[66]; // @[BOOTH_gen.scala 29:20]
  assign RS_66_io_x_sub = io_x[65]; // @[BOOTH_gen.scala 30:24]
  assign RS_67_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_67_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_67_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_67_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_67_io_x = io_x[67]; // @[BOOTH_gen.scala 29:20]
  assign RS_67_io_x_sub = io_x[66]; // @[BOOTH_gen.scala 30:24]
  assign RS_68_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_68_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_68_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_68_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_68_io_x = io_x[68]; // @[BOOTH_gen.scala 29:20]
  assign RS_68_io_x_sub = io_x[67]; // @[BOOTH_gen.scala 30:24]
  assign RS_69_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_69_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_69_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_69_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_69_io_x = io_x[69]; // @[BOOTH_gen.scala 29:20]
  assign RS_69_io_x_sub = io_x[68]; // @[BOOTH_gen.scala 30:24]
  assign RS_70_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_70_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_70_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_70_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_70_io_x = io_x[70]; // @[BOOTH_gen.scala 29:20]
  assign RS_70_io_x_sub = io_x[69]; // @[BOOTH_gen.scala 30:24]
  assign RS_71_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_71_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_71_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_71_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_71_io_x = io_x[71]; // @[BOOTH_gen.scala 29:20]
  assign RS_71_io_x_sub = io_x[70]; // @[BOOTH_gen.scala 30:24]
  assign RS_72_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_72_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_72_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_72_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_72_io_x = io_x[72]; // @[BOOTH_gen.scala 29:20]
  assign RS_72_io_x_sub = io_x[71]; // @[BOOTH_gen.scala 30:24]
  assign RS_73_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_73_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_73_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_73_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_73_io_x = io_x[73]; // @[BOOTH_gen.scala 29:20]
  assign RS_73_io_x_sub = io_x[72]; // @[BOOTH_gen.scala 30:24]
  assign RS_74_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_74_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_74_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_74_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_74_io_x = io_x[74]; // @[BOOTH_gen.scala 29:20]
  assign RS_74_io_x_sub = io_x[73]; // @[BOOTH_gen.scala 30:24]
  assign RS_75_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_75_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_75_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_75_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_75_io_x = io_x[75]; // @[BOOTH_gen.scala 29:20]
  assign RS_75_io_x_sub = io_x[74]; // @[BOOTH_gen.scala 30:24]
  assign RS_76_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_76_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_76_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_76_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_76_io_x = io_x[76]; // @[BOOTH_gen.scala 29:20]
  assign RS_76_io_x_sub = io_x[75]; // @[BOOTH_gen.scala 30:24]
  assign RS_77_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_77_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_77_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_77_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_77_io_x = io_x[77]; // @[BOOTH_gen.scala 29:20]
  assign RS_77_io_x_sub = io_x[76]; // @[BOOTH_gen.scala 30:24]
  assign RS_78_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_78_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_78_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_78_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_78_io_x = io_x[78]; // @[BOOTH_gen.scala 29:20]
  assign RS_78_io_x_sub = io_x[77]; // @[BOOTH_gen.scala 30:24]
  assign RS_79_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_79_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_79_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_79_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_79_io_x = io_x[79]; // @[BOOTH_gen.scala 29:20]
  assign RS_79_io_x_sub = io_x[78]; // @[BOOTH_gen.scala 30:24]
  assign RS_80_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_80_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_80_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_80_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_80_io_x = io_x[80]; // @[BOOTH_gen.scala 29:20]
  assign RS_80_io_x_sub = io_x[79]; // @[BOOTH_gen.scala 30:24]
  assign RS_81_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_81_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_81_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_81_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_81_io_x = io_x[81]; // @[BOOTH_gen.scala 29:20]
  assign RS_81_io_x_sub = io_x[80]; // @[BOOTH_gen.scala 30:24]
  assign RS_82_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_82_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_82_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_82_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_82_io_x = io_x[82]; // @[BOOTH_gen.scala 29:20]
  assign RS_82_io_x_sub = io_x[81]; // @[BOOTH_gen.scala 30:24]
  assign RS_83_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_83_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_83_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_83_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_83_io_x = io_x[83]; // @[BOOTH_gen.scala 29:20]
  assign RS_83_io_x_sub = io_x[82]; // @[BOOTH_gen.scala 30:24]
  assign RS_84_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_84_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_84_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_84_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_84_io_x = io_x[84]; // @[BOOTH_gen.scala 29:20]
  assign RS_84_io_x_sub = io_x[83]; // @[BOOTH_gen.scala 30:24]
  assign RS_85_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_85_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_85_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_85_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_85_io_x = io_x[85]; // @[BOOTH_gen.scala 29:20]
  assign RS_85_io_x_sub = io_x[84]; // @[BOOTH_gen.scala 30:24]
  assign RS_86_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_86_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_86_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_86_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_86_io_x = io_x[86]; // @[BOOTH_gen.scala 29:20]
  assign RS_86_io_x_sub = io_x[85]; // @[BOOTH_gen.scala 30:24]
  assign RS_87_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_87_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_87_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_87_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_87_io_x = io_x[87]; // @[BOOTH_gen.scala 29:20]
  assign RS_87_io_x_sub = io_x[86]; // @[BOOTH_gen.scala 30:24]
  assign RS_88_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_88_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_88_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_88_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_88_io_x = io_x[88]; // @[BOOTH_gen.scala 29:20]
  assign RS_88_io_x_sub = io_x[87]; // @[BOOTH_gen.scala 30:24]
  assign RS_89_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_89_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_89_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_89_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_89_io_x = io_x[89]; // @[BOOTH_gen.scala 29:20]
  assign RS_89_io_x_sub = io_x[88]; // @[BOOTH_gen.scala 30:24]
  assign RS_90_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_90_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_90_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_90_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_90_io_x = io_x[90]; // @[BOOTH_gen.scala 29:20]
  assign RS_90_io_x_sub = io_x[89]; // @[BOOTH_gen.scala 30:24]
  assign RS_91_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_91_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_91_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_91_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_91_io_x = io_x[91]; // @[BOOTH_gen.scala 29:20]
  assign RS_91_io_x_sub = io_x[90]; // @[BOOTH_gen.scala 30:24]
  assign RS_92_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_92_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_92_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_92_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_92_io_x = io_x[92]; // @[BOOTH_gen.scala 29:20]
  assign RS_92_io_x_sub = io_x[91]; // @[BOOTH_gen.scala 30:24]
  assign RS_93_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_93_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_93_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_93_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_93_io_x = io_x[93]; // @[BOOTH_gen.scala 29:20]
  assign RS_93_io_x_sub = io_x[92]; // @[BOOTH_gen.scala 30:24]
  assign RS_94_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_94_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_94_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_94_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_94_io_x = io_x[94]; // @[BOOTH_gen.scala 29:20]
  assign RS_94_io_x_sub = io_x[93]; // @[BOOTH_gen.scala 30:24]
  assign RS_95_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_95_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_95_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_95_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_95_io_x = io_x[95]; // @[BOOTH_gen.scala 29:20]
  assign RS_95_io_x_sub = io_x[94]; // @[BOOTH_gen.scala 30:24]
  assign RS_96_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_96_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_96_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_96_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_96_io_x = io_x[96]; // @[BOOTH_gen.scala 29:20]
  assign RS_96_io_x_sub = io_x[95]; // @[BOOTH_gen.scala 30:24]
  assign RS_97_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_97_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_97_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_97_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_97_io_x = io_x[97]; // @[BOOTH_gen.scala 29:20]
  assign RS_97_io_x_sub = io_x[96]; // @[BOOTH_gen.scala 30:24]
  assign RS_98_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_98_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_98_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_98_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_98_io_x = io_x[98]; // @[BOOTH_gen.scala 29:20]
  assign RS_98_io_x_sub = io_x[97]; // @[BOOTH_gen.scala 30:24]
  assign RS_99_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_99_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_99_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_99_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_99_io_x = io_x[99]; // @[BOOTH_gen.scala 29:20]
  assign RS_99_io_x_sub = io_x[98]; // @[BOOTH_gen.scala 30:24]
  assign RS_100_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_100_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_100_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_100_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_100_io_x = io_x[100]; // @[BOOTH_gen.scala 29:20]
  assign RS_100_io_x_sub = io_x[99]; // @[BOOTH_gen.scala 30:24]
  assign RS_101_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_101_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_101_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_101_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_101_io_x = io_x[101]; // @[BOOTH_gen.scala 29:20]
  assign RS_101_io_x_sub = io_x[100]; // @[BOOTH_gen.scala 30:24]
  assign RS_102_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_102_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_102_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_102_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_102_io_x = io_x[102]; // @[BOOTH_gen.scala 29:20]
  assign RS_102_io_x_sub = io_x[101]; // @[BOOTH_gen.scala 30:24]
  assign RS_103_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_103_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_103_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_103_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_103_io_x = io_x[103]; // @[BOOTH_gen.scala 29:20]
  assign RS_103_io_x_sub = io_x[102]; // @[BOOTH_gen.scala 30:24]
  assign RS_104_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_104_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_104_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_104_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_104_io_x = io_x[104]; // @[BOOTH_gen.scala 29:20]
  assign RS_104_io_x_sub = io_x[103]; // @[BOOTH_gen.scala 30:24]
  assign RS_105_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_105_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_105_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_105_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_105_io_x = io_x[105]; // @[BOOTH_gen.scala 29:20]
  assign RS_105_io_x_sub = io_x[104]; // @[BOOTH_gen.scala 30:24]
  assign RS_106_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_106_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_106_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_106_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_106_io_x = io_x[106]; // @[BOOTH_gen.scala 29:20]
  assign RS_106_io_x_sub = io_x[105]; // @[BOOTH_gen.scala 30:24]
  assign RS_107_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_107_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_107_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_107_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_107_io_x = io_x[107]; // @[BOOTH_gen.scala 29:20]
  assign RS_107_io_x_sub = io_x[106]; // @[BOOTH_gen.scala 30:24]
  assign RS_108_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_108_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_108_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_108_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_108_io_x = io_x[108]; // @[BOOTH_gen.scala 29:20]
  assign RS_108_io_x_sub = io_x[107]; // @[BOOTH_gen.scala 30:24]
  assign RS_109_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_109_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_109_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_109_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_109_io_x = io_x[109]; // @[BOOTH_gen.scala 29:20]
  assign RS_109_io_x_sub = io_x[108]; // @[BOOTH_gen.scala 30:24]
  assign RS_110_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_110_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_110_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_110_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_110_io_x = io_x[110]; // @[BOOTH_gen.scala 29:20]
  assign RS_110_io_x_sub = io_x[109]; // @[BOOTH_gen.scala 30:24]
  assign RS_111_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_111_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_111_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_111_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_111_io_x = io_x[111]; // @[BOOTH_gen.scala 29:20]
  assign RS_111_io_x_sub = io_x[110]; // @[BOOTH_gen.scala 30:24]
  assign RS_112_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_112_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_112_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_112_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_112_io_x = io_x[112]; // @[BOOTH_gen.scala 29:20]
  assign RS_112_io_x_sub = io_x[111]; // @[BOOTH_gen.scala 30:24]
  assign RS_113_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_113_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_113_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_113_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_113_io_x = io_x[113]; // @[BOOTH_gen.scala 29:20]
  assign RS_113_io_x_sub = io_x[112]; // @[BOOTH_gen.scala 30:24]
  assign RS_114_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_114_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_114_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_114_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_114_io_x = io_x[114]; // @[BOOTH_gen.scala 29:20]
  assign RS_114_io_x_sub = io_x[113]; // @[BOOTH_gen.scala 30:24]
  assign RS_115_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_115_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_115_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_115_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_115_io_x = io_x[115]; // @[BOOTH_gen.scala 29:20]
  assign RS_115_io_x_sub = io_x[114]; // @[BOOTH_gen.scala 30:24]
  assign RS_116_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_116_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_116_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_116_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_116_io_x = io_x[116]; // @[BOOTH_gen.scala 29:20]
  assign RS_116_io_x_sub = io_x[115]; // @[BOOTH_gen.scala 30:24]
  assign RS_117_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_117_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_117_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_117_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_117_io_x = io_x[117]; // @[BOOTH_gen.scala 29:20]
  assign RS_117_io_x_sub = io_x[116]; // @[BOOTH_gen.scala 30:24]
  assign RS_118_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_118_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_118_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_118_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_118_io_x = io_x[118]; // @[BOOTH_gen.scala 29:20]
  assign RS_118_io_x_sub = io_x[117]; // @[BOOTH_gen.scala 30:24]
  assign RS_119_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_119_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_119_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_119_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_119_io_x = io_x[119]; // @[BOOTH_gen.scala 29:20]
  assign RS_119_io_x_sub = io_x[118]; // @[BOOTH_gen.scala 30:24]
  assign RS_120_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_120_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_120_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_120_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_120_io_x = io_x[120]; // @[BOOTH_gen.scala 29:20]
  assign RS_120_io_x_sub = io_x[119]; // @[BOOTH_gen.scala 30:24]
  assign RS_121_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_121_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_121_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_121_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_121_io_x = io_x[121]; // @[BOOTH_gen.scala 29:20]
  assign RS_121_io_x_sub = io_x[120]; // @[BOOTH_gen.scala 30:24]
  assign RS_122_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_122_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_122_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_122_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_122_io_x = io_x[122]; // @[BOOTH_gen.scala 29:20]
  assign RS_122_io_x_sub = io_x[121]; // @[BOOTH_gen.scala 30:24]
  assign RS_123_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_123_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_123_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_123_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_123_io_x = io_x[123]; // @[BOOTH_gen.scala 29:20]
  assign RS_123_io_x_sub = io_x[122]; // @[BOOTH_gen.scala 30:24]
  assign RS_124_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_124_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_124_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_124_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_124_io_x = io_x[124]; // @[BOOTH_gen.scala 29:20]
  assign RS_124_io_x_sub = io_x[123]; // @[BOOTH_gen.scala 30:24]
  assign RS_125_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_125_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_125_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_125_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_125_io_x = io_x[125]; // @[BOOTH_gen.scala 29:20]
  assign RS_125_io_x_sub = io_x[124]; // @[BOOTH_gen.scala 30:24]
  assign RS_126_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_126_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_126_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_126_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_126_io_x = io_x[126]; // @[BOOTH_gen.scala 29:20]
  assign RS_126_io_x_sub = io_x[125]; // @[BOOTH_gen.scala 30:24]
  assign RS_127_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_127_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_127_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_127_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_127_io_x = io_x[127]; // @[BOOTH_gen.scala 29:20]
  assign RS_127_io_x_sub = io_x[126]; // @[BOOTH_gen.scala 30:24]
  assign RS_128_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_128_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_128_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_128_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_128_io_x = io_x[128]; // @[BOOTH_gen.scala 29:20]
  assign RS_128_io_x_sub = io_x[127]; // @[BOOTH_gen.scala 30:24]
  assign RS_129_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_129_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_129_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_129_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_129_io_x = io_x[129]; // @[BOOTH_gen.scala 29:20]
  assign RS_129_io_x_sub = io_x[128]; // @[BOOTH_gen.scala 30:24]
  assign RS_130_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_130_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_130_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_130_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_130_io_x = io_x[130]; // @[BOOTH_gen.scala 29:20]
  assign RS_130_io_x_sub = io_x[129]; // @[BOOTH_gen.scala 30:24]
  assign RS_131_io_sel_negative = BOOTH_S_io_sel_negative; // @[BOOTH_gen.scala 16:20 31:27]
  assign RS_131_io_sel_positive = BOOTH_S_io_sel_positive; // @[BOOTH_gen.scala 16:20 32:27]
  assign RS_131_io_sel_double_negative = BOOTH_S_io_sel_double_negative; // @[BOOTH_gen.scala 16:20 33:34]
  assign RS_131_io_sel_double_positive = BOOTH_S_io_sel_double_positive; // @[BOOTH_gen.scala 16:20 34:34]
  assign RS_131_io_x = io_x[131]; // @[BOOTH_gen.scala 29:20]
  assign RS_131_io_x_sub = io_x[130]; // @[BOOTH_gen.scala 30:24]
  assign BOOTH_S_io_src = io_y; // @[BOOTH_gen.scala 19:11]
endmodule
module mul(
  input         clock,
  input         reset,
  input         io_mul_valid,
  input  [63:0] io_multiplicand,
  input  [63:0] io_multiplier,
  output        io_out_valid,
  output [63:0] io_result_lo
);
`ifdef RANDOMIZE_REG_INIT
  reg [159:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [131:0] BOOTH_gen_io_x; // @[mul.scala 101:18]
  wire [2:0] BOOTH_gen_io_y; // @[mul.scala 101:18]
  wire [131:0] BOOTH_gen_io_out; // @[mul.scala 101:18]
  wire  BOOTH_gen_io_cout; // @[mul.scala 101:18]
  wire [65:0] multiplier = {io_multiplier[63],io_multiplier,1'h0}; // @[Cat.scala 31:58]
  wire [65:0] multiplicand = {io_multiplicand[63],io_multiplicand,1'h0}; // @[Cat.scala 31:58]
  reg [131:0] multiplicand_reg; // @[mul.scala 75:33]
  reg [65:0] multiplier_reg; // @[mul.scala 76:33]
  reg [131:0] result; // @[mul.scala 77:33]
  reg  start; // @[mul.scala 78:33]
  wire  _GEN_1 = io_mul_valid | start; // @[mul.scala 81:22 83:18 78:33]
  wire  _multiplier_reg_T_1 = ~start & io_mul_valid; // @[mul.scala 98:45]
  wire [133:0] _multiplicand_reg_T_2 = {multiplicand_reg, 2'h0}; // @[mul.scala 99:93]
  wire [133:0] _multiplicand_reg_T_3 = _multiplier_reg_T_1 ? {{68'd0}, multiplicand} : _multiplicand_reg_T_2; // @[mul.scala 99:26]
  wire [131:0] _result_T_2 = result + BOOTH_gen_io_out; // @[mul.scala 105:42]
  wire [131:0] _GEN_0 = {{131'd0}, BOOTH_gen_io_cout}; // @[mul.scala 105:51]
  wire [131:0] _result_T_4 = _result_T_2 + _GEN_0; // @[mul.scala 105:51]
  wire  result_sign = io_multiplier[63] ^ io_multiplicand[63]; // @[mul.scala 108:30]
  wire [133:0] _GEN_6 = reset ? 134'h0 : _multiplicand_reg_T_3; // @[mul.scala 75:{33,33} 99:20]
  BOOTH_gen BOOTH_gen ( // @[mul.scala 101:18]
    .io_x(BOOTH_gen_io_x),
    .io_y(BOOTH_gen_io_y),
    .io_out(BOOTH_gen_io_out),
    .io_cout(BOOTH_gen_io_cout)
  );
  assign io_out_valid = multiplier_reg == 66'h0 & start; // @[mul.scala 87:31]
  assign io_result_lo = {result_sign,result[63:1]}; // @[Cat.scala 31:58]
  assign BOOTH_gen_io_x = multiplicand_reg; // @[mul.scala 103:8]
  assign BOOTH_gen_io_y = multiplier_reg[2:0]; // @[mul.scala 102:25]
  always @(posedge clock) begin
    multiplicand_reg <= _GEN_6[131:0]; // @[mul.scala 75:{33,33} 99:20]
    if (reset) begin // @[mul.scala 76:33]
      multiplier_reg <= 66'h0; // @[mul.scala 76:33]
    end else if (~start & io_mul_valid) begin // @[mul.scala 98:26]
      multiplier_reg <= multiplier;
    end else begin
      multiplier_reg <= {{2'd0}, multiplier_reg[65:2]};
    end
    if (reset) begin // @[mul.scala 77:33]
      result <= 132'h0; // @[mul.scala 77:33]
    end else if (io_out_valid) begin // @[mul.scala 113:21]
      result <= 132'h0; // @[mul.scala 114:12]
    end else if (start) begin // @[mul.scala 105:16]
      result <= _result_T_4;
    end
    if (reset) begin // @[mul.scala 78:33]
      start <= 1'h0; // @[mul.scala 78:33]
    end else if (multiplier_reg == 66'h0 & start) begin // @[mul.scala 87:52]
      start <= 1'h0; // @[mul.scala 90:18]
    end else begin
      start <= _GEN_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {5{`RANDOM}};
  multiplicand_reg = _RAND_0[131:0];
  _RAND_1 = {3{`RANDOM}};
  multiplier_reg = _RAND_1[65:0];
  _RAND_2 = {5{`RANDOM}};
  result = _RAND_2[131:0];
  _RAND_3 = {1{`RANDOM}};
  start = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module mul_1(
  input         clock,
  input         reset,
  input         io_mul_valid,
  input  [31:0] io_multiplicand,
  input  [31:0] io_multiplier,
  output        io_out_valid,
  output [31:0] io_result_lo
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [131:0] BOOTH_gen_io_x; // @[mul.scala 101:18]
  wire [2:0] BOOTH_gen_io_y; // @[mul.scala 101:18]
  wire [131:0] BOOTH_gen_io_out; // @[mul.scala 101:18]
  wire  BOOTH_gen_io_cout; // @[mul.scala 101:18]
  wire [33:0] multiplier = {1'h0,io_multiplier,1'h0}; // @[Cat.scala 31:58]
  wire [33:0] multiplicand = {1'h0,io_multiplicand,1'h0}; // @[Cat.scala 31:58]
  reg [67:0] multiplicand_reg; // @[mul.scala 75:33]
  reg [33:0] multiplier_reg; // @[mul.scala 76:33]
  reg [67:0] result; // @[mul.scala 77:33]
  reg  start; // @[mul.scala 78:33]
  wire  _GEN_1 = io_mul_valid | start; // @[mul.scala 81:22 83:18 78:33]
  wire  _multiplier_reg_T_1 = ~start & io_mul_valid; // @[mul.scala 98:45]
  wire [69:0] _multiplicand_reg_T_2 = {multiplicand_reg, 2'h0}; // @[mul.scala 99:93]
  wire [69:0] _multiplicand_reg_T_3 = _multiplier_reg_T_1 ? {{36'd0}, multiplicand} : _multiplicand_reg_T_2; // @[mul.scala 99:26]
  wire [131:0] _GEN_0 = {{64'd0}, result}; // @[mul.scala 105:42]
  wire [131:0] _result_T_2 = _GEN_0 + BOOTH_gen_io_out; // @[mul.scala 105:42]
  wire [131:0] _GEN_6 = {{131'd0}, BOOTH_gen_io_cout}; // @[mul.scala 105:51]
  wire [131:0] _result_T_4 = _result_T_2 + _GEN_6; // @[mul.scala 105:51]
  wire [131:0] _result_T_5 = start ? _result_T_4 : {{64'd0}, result}; // @[mul.scala 105:16]
  wire  result_sign = io_multiplier[31] ^ io_multiplicand[31]; // @[mul.scala 108:30]
  wire [131:0] _GEN_5 = io_out_valid ? 132'h0 : _result_T_5; // @[mul.scala 105:10 113:21 114:12]
  wire [69:0] _GEN_7 = reset ? 70'h0 : _multiplicand_reg_T_3; // @[mul.scala 75:{33,33} 99:20]
  wire [131:0] _GEN_8 = reset ? 132'h0 : _GEN_5; // @[mul.scala 77:{33,33}]
  BOOTH_gen BOOTH_gen ( // @[mul.scala 101:18]
    .io_x(BOOTH_gen_io_x),
    .io_y(BOOTH_gen_io_y),
    .io_out(BOOTH_gen_io_out),
    .io_cout(BOOTH_gen_io_cout)
  );
  assign io_out_valid = multiplier_reg == 34'h0 & start; // @[mul.scala 87:31]
  assign io_result_lo = {result_sign,result[31:1]}; // @[Cat.scala 31:58]
  assign BOOTH_gen_io_x = {{64'd0}, multiplicand_reg}; // @[mul.scala 103:8]
  assign BOOTH_gen_io_y = multiplier_reg[2:0]; // @[mul.scala 102:25]
  always @(posedge clock) begin
    multiplicand_reg <= _GEN_7[67:0]; // @[mul.scala 75:{33,33} 99:20]
    if (reset) begin // @[mul.scala 76:33]
      multiplier_reg <= 34'h0; // @[mul.scala 76:33]
    end else if (~start & io_mul_valid) begin // @[mul.scala 98:26]
      multiplier_reg <= multiplier;
    end else begin
      multiplier_reg <= {{2'd0}, multiplier_reg[33:2]};
    end
    result <= _GEN_8[67:0]; // @[mul.scala 77:{33,33}]
    if (reset) begin // @[mul.scala 78:33]
      start <= 1'h0; // @[mul.scala 78:33]
    end else if (multiplier_reg == 34'h0 & start) begin // @[mul.scala 87:52]
      start <= 1'h0; // @[mul.scala 90:18]
    end else begin
      start <= _GEN_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  multiplicand_reg = _RAND_0[67:0];
  _RAND_1 = {2{`RANDOM}};
  multiplier_reg = _RAND_1[33:0];
  _RAND_2 = {3{`RANDOM}};
  result = _RAND_2[67:0];
  _RAND_3 = {1{`RANDOM}};
  start = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module div(
  input         clock,
  input         reset,
  input  [63:0] io_dividend,
  input  [63:0] io_divisor,
  input         io_div_valid,
  input         io_div_signed,
  output        io_out_valid,
  output [63:0] io_quotient,
  output [63:0] io_remainder
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [127:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] dividend_reg; // @[div.scala 21:25]
  reg [63:0] divisor_reg; // @[div.scala 22:25]
  reg  start; // @[div.scala 23:25]
  reg [7:0] delay; // @[div.scala 25:24]
  reg [1:0] clear; // @[div.scala 27:24]
  wire  _dividend_T_1 = io_div_signed & io_dividend[63]; // @[div.scala 31:34]
  wire [63:0] _dividend_T_3 = ~io_dividend; // @[div.scala 31:66]
  wire [63:0] _dividend_T_5 = _dividend_T_3 + 64'h1; // @[div.scala 31:80]
  wire [63:0] _divisor_T_3 = ~io_divisor; // @[div.scala 32:65]
  wire [63:0] _divisor_T_5 = _divisor_T_3 + 64'h1; // @[div.scala 32:78]
  reg  quotient_sign; // @[div.scala 42:31]
  reg  remainder_sign; // @[div.scala 43:31]
  reg [127:0] A; // @[div.scala 48:18]
  reg [63:0] B; // @[div.scala 49:18]
  reg [63:0] S; // @[div.scala 51:18]
  reg [7:0] cnt; // @[div.scala 52:20]
  wire [127:0] _A_T = {64'h0,dividend_reg}; // @[Cat.scala 31:58]
  wire  _T_1 = ~io_out_valid; // @[div.scala 58:23]
  wire [7:0] _delay_T_1 = delay + 8'h1; // @[div.scala 59:20]
  wire [64:0] _S_tmp_T_1 = {1'h0,B}; // @[Cat.scala 31:58]
  wire  _S_tmp_T_2 = A[127:63] >= _S_tmp_T_1; // @[div.scala 61:42]
  wire  _GEN_3 = 6'h0 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_4 = 6'h1 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_5 = 6'h2 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_6 = 6'h3 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_7 = 6'h4 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_8 = 6'h5 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_9 = 6'h6 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_10 = 6'h7 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_11 = 6'h8 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_12 = 6'h9 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_13 = 6'ha == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_14 = 6'hb == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_15 = 6'hc == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_16 = 6'hd == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_17 = 6'he == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_18 = 6'hf == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_19 = 6'h10 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_20 = 6'h11 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_21 = 6'h12 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_22 = 6'h13 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_23 = 6'h14 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_24 = 6'h15 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_25 = 6'h16 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_26 = 6'h17 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_27 = 6'h18 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_28 = 6'h19 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_29 = 6'h1a == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_30 = 6'h1b == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_31 = 6'h1c == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_32 = 6'h1d == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_33 = 6'h1e == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_34 = 6'h1f == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_35 = 6'h20 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_36 = 6'h21 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_37 = 6'h22 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_38 = 6'h23 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_39 = 6'h24 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_40 = 6'h25 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_41 = 6'h26 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_42 = 6'h27 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_43 = 6'h28 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_44 = 6'h29 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_45 = 6'h2a == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_46 = 6'h2b == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_47 = 6'h2c == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_48 = 6'h2d == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_49 = 6'h2e == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_50 = 6'h2f == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_51 = 6'h30 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_52 = 6'h31 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_53 = 6'h32 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_54 = 6'h33 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_55 = 6'h34 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_56 = 6'h35 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_57 = 6'h36 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_58 = 6'h37 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_59 = 6'h38 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_60 = 6'h39 == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_61 = 6'h3a == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_62 = 6'h3b == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_63 = 6'h3c == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_64 = 6'h3d == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_65 = 6'h3e == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_66 = 6'h3f == cnt[5:0] & A[127:63] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire [127:0] _A_T_5 = {65'h0,A[62:0]}; // @[Cat.scala 31:58]
  wire [64:0] _A_T_9 = A[127:63] - _S_tmp_T_1; // @[div.scala 62:106]
  wire [127:0] _A_T_10 = {_A_T_9, 63'h0}; // @[div.scala 62:121]
  wire [127:0] _A_T_11 = _A_T_5 | _A_T_10; // @[div.scala 62:84]
  wire [127:0] _A_T_12 = _S_tmp_T_2 ? _A_T_11 : A; // @[div.scala 62:14]
  wire [128:0] _A_T_13 = {_A_T_12, 1'h0}; // @[div.scala 62:137]
  wire [7:0] _cnt_T_1 = cnt + 8'h1; // @[div.scala 63:16]
  wire  _GEN_129 = delay >= 8'h2 & _T_1 & _GEN_65; // @[div.scala 50:22 60:44]
  wire  S_tmp_62 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_129; // @[div.scala 50:22 58:46]
  wire  _GEN_130 = delay >= 8'h2 & _T_1 & _GEN_66; // @[div.scala 50:22 60:44]
  wire  S_tmp_63 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_130; // @[div.scala 50:22 58:46]
  wire  _GEN_127 = delay >= 8'h2 & _T_1 & _GEN_63; // @[div.scala 50:22 60:44]
  wire  S_tmp_60 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_127; // @[div.scala 50:22 58:46]
  wire  _GEN_128 = delay >= 8'h2 & _T_1 & _GEN_64; // @[div.scala 50:22 60:44]
  wire  S_tmp_61 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_128; // @[div.scala 50:22 58:46]
  wire  _GEN_125 = delay >= 8'h2 & _T_1 & _GEN_61; // @[div.scala 50:22 60:44]
  wire  S_tmp_58 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_125; // @[div.scala 50:22 58:46]
  wire  _GEN_126 = delay >= 8'h2 & _T_1 & _GEN_62; // @[div.scala 50:22 60:44]
  wire  S_tmp_59 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_126; // @[div.scala 50:22 58:46]
  wire  _GEN_123 = delay >= 8'h2 & _T_1 & _GEN_59; // @[div.scala 50:22 60:44]
  wire  S_tmp_56 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_123; // @[div.scala 50:22 58:46]
  wire  _GEN_124 = delay >= 8'h2 & _T_1 & _GEN_60; // @[div.scala 50:22 60:44]
  wire  S_tmp_57 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_124; // @[div.scala 50:22 58:46]
  wire [7:0] S_lo_lo_lo = {S_tmp_56,S_tmp_57,S_tmp_58,S_tmp_59,S_tmp_60,S_tmp_61,S_tmp_62,S_tmp_63}; // @[Cat.scala 31:58]
  wire  _GEN_121 = delay >= 8'h2 & _T_1 & _GEN_57; // @[div.scala 50:22 60:44]
  wire  S_tmp_54 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_121; // @[div.scala 50:22 58:46]
  wire  _GEN_122 = delay >= 8'h2 & _T_1 & _GEN_58; // @[div.scala 50:22 60:44]
  wire  S_tmp_55 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_122; // @[div.scala 50:22 58:46]
  wire  _GEN_119 = delay >= 8'h2 & _T_1 & _GEN_55; // @[div.scala 50:22 60:44]
  wire  S_tmp_52 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_119; // @[div.scala 50:22 58:46]
  wire  _GEN_120 = delay >= 8'h2 & _T_1 & _GEN_56; // @[div.scala 50:22 60:44]
  wire  S_tmp_53 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_120; // @[div.scala 50:22 58:46]
  wire  _GEN_117 = delay >= 8'h2 & _T_1 & _GEN_53; // @[div.scala 50:22 60:44]
  wire  S_tmp_50 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_117; // @[div.scala 50:22 58:46]
  wire  _GEN_118 = delay >= 8'h2 & _T_1 & _GEN_54; // @[div.scala 50:22 60:44]
  wire  S_tmp_51 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_118; // @[div.scala 50:22 58:46]
  wire  _GEN_115 = delay >= 8'h2 & _T_1 & _GEN_51; // @[div.scala 50:22 60:44]
  wire  S_tmp_48 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_115; // @[div.scala 50:22 58:46]
  wire  _GEN_116 = delay >= 8'h2 & _T_1 & _GEN_52; // @[div.scala 50:22 60:44]
  wire  S_tmp_49 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_116; // @[div.scala 50:22 58:46]
  wire [15:0] S_lo_lo = {S_tmp_48,S_tmp_49,S_tmp_50,S_tmp_51,S_tmp_52,S_tmp_53,S_tmp_54,S_tmp_55,S_lo_lo_lo}; // @[Cat.scala 31:58]
  wire  _GEN_113 = delay >= 8'h2 & _T_1 & _GEN_49; // @[div.scala 50:22 60:44]
  wire  S_tmp_46 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_113; // @[div.scala 50:22 58:46]
  wire  _GEN_114 = delay >= 8'h2 & _T_1 & _GEN_50; // @[div.scala 50:22 60:44]
  wire  S_tmp_47 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_114; // @[div.scala 50:22 58:46]
  wire  _GEN_111 = delay >= 8'h2 & _T_1 & _GEN_47; // @[div.scala 50:22 60:44]
  wire  S_tmp_44 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_111; // @[div.scala 50:22 58:46]
  wire  _GEN_112 = delay >= 8'h2 & _T_1 & _GEN_48; // @[div.scala 50:22 60:44]
  wire  S_tmp_45 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_112; // @[div.scala 50:22 58:46]
  wire  _GEN_109 = delay >= 8'h2 & _T_1 & _GEN_45; // @[div.scala 50:22 60:44]
  wire  S_tmp_42 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_109; // @[div.scala 50:22 58:46]
  wire  _GEN_110 = delay >= 8'h2 & _T_1 & _GEN_46; // @[div.scala 50:22 60:44]
  wire  S_tmp_43 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_110; // @[div.scala 50:22 58:46]
  wire  _GEN_107 = delay >= 8'h2 & _T_1 & _GEN_43; // @[div.scala 50:22 60:44]
  wire  S_tmp_40 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_107; // @[div.scala 50:22 58:46]
  wire  _GEN_108 = delay >= 8'h2 & _T_1 & _GEN_44; // @[div.scala 50:22 60:44]
  wire  S_tmp_41 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_108; // @[div.scala 50:22 58:46]
  wire [7:0] S_lo_hi_lo = {S_tmp_40,S_tmp_41,S_tmp_42,S_tmp_43,S_tmp_44,S_tmp_45,S_tmp_46,S_tmp_47}; // @[Cat.scala 31:58]
  wire  _GEN_105 = delay >= 8'h2 & _T_1 & _GEN_41; // @[div.scala 50:22 60:44]
  wire  S_tmp_38 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_105; // @[div.scala 50:22 58:46]
  wire  _GEN_106 = delay >= 8'h2 & _T_1 & _GEN_42; // @[div.scala 50:22 60:44]
  wire  S_tmp_39 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_106; // @[div.scala 50:22 58:46]
  wire  _GEN_103 = delay >= 8'h2 & _T_1 & _GEN_39; // @[div.scala 50:22 60:44]
  wire  S_tmp_36 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_103; // @[div.scala 50:22 58:46]
  wire  _GEN_104 = delay >= 8'h2 & _T_1 & _GEN_40; // @[div.scala 50:22 60:44]
  wire  S_tmp_37 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_104; // @[div.scala 50:22 58:46]
  wire  _GEN_101 = delay >= 8'h2 & _T_1 & _GEN_37; // @[div.scala 50:22 60:44]
  wire  S_tmp_34 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_101; // @[div.scala 50:22 58:46]
  wire  _GEN_102 = delay >= 8'h2 & _T_1 & _GEN_38; // @[div.scala 50:22 60:44]
  wire  S_tmp_35 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_102; // @[div.scala 50:22 58:46]
  wire  _GEN_99 = delay >= 8'h2 & _T_1 & _GEN_35; // @[div.scala 50:22 60:44]
  wire  S_tmp_32 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_99; // @[div.scala 50:22 58:46]
  wire  _GEN_100 = delay >= 8'h2 & _T_1 & _GEN_36; // @[div.scala 50:22 60:44]
  wire  S_tmp_33 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_100; // @[div.scala 50:22 58:46]
  wire [31:0] S_lo = {S_tmp_32,S_tmp_33,S_tmp_34,S_tmp_35,S_tmp_36,S_tmp_37,S_tmp_38,S_tmp_39,S_lo_hi_lo,S_lo_lo}; // @[Cat.scala 31:58]
  wire  _GEN_97 = delay >= 8'h2 & _T_1 & _GEN_33; // @[div.scala 50:22 60:44]
  wire  S_tmp_30 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_97; // @[div.scala 50:22 58:46]
  wire  _GEN_98 = delay >= 8'h2 & _T_1 & _GEN_34; // @[div.scala 50:22 60:44]
  wire  S_tmp_31 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_98; // @[div.scala 50:22 58:46]
  wire  _GEN_95 = delay >= 8'h2 & _T_1 & _GEN_31; // @[div.scala 50:22 60:44]
  wire  S_tmp_28 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_95; // @[div.scala 50:22 58:46]
  wire  _GEN_96 = delay >= 8'h2 & _T_1 & _GEN_32; // @[div.scala 50:22 60:44]
  wire  S_tmp_29 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_96; // @[div.scala 50:22 58:46]
  wire  _GEN_93 = delay >= 8'h2 & _T_1 & _GEN_29; // @[div.scala 50:22 60:44]
  wire  S_tmp_26 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_93; // @[div.scala 50:22 58:46]
  wire  _GEN_94 = delay >= 8'h2 & _T_1 & _GEN_30; // @[div.scala 50:22 60:44]
  wire  S_tmp_27 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_94; // @[div.scala 50:22 58:46]
  wire  _GEN_91 = delay >= 8'h2 & _T_1 & _GEN_27; // @[div.scala 50:22 60:44]
  wire  S_tmp_24 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_91; // @[div.scala 50:22 58:46]
  wire  _GEN_92 = delay >= 8'h2 & _T_1 & _GEN_28; // @[div.scala 50:22 60:44]
  wire  S_tmp_25 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_92; // @[div.scala 50:22 58:46]
  wire [7:0] S_hi_lo_lo = {S_tmp_24,S_tmp_25,S_tmp_26,S_tmp_27,S_tmp_28,S_tmp_29,S_tmp_30,S_tmp_31}; // @[Cat.scala 31:58]
  wire  _GEN_89 = delay >= 8'h2 & _T_1 & _GEN_25; // @[div.scala 50:22 60:44]
  wire  S_tmp_22 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_89; // @[div.scala 50:22 58:46]
  wire  _GEN_90 = delay >= 8'h2 & _T_1 & _GEN_26; // @[div.scala 50:22 60:44]
  wire  S_tmp_23 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_90; // @[div.scala 50:22 58:46]
  wire  _GEN_87 = delay >= 8'h2 & _T_1 & _GEN_23; // @[div.scala 50:22 60:44]
  wire  S_tmp_20 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_87; // @[div.scala 50:22 58:46]
  wire  _GEN_88 = delay >= 8'h2 & _T_1 & _GEN_24; // @[div.scala 50:22 60:44]
  wire  S_tmp_21 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_88; // @[div.scala 50:22 58:46]
  wire  _GEN_85 = delay >= 8'h2 & _T_1 & _GEN_21; // @[div.scala 50:22 60:44]
  wire  S_tmp_18 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_85; // @[div.scala 50:22 58:46]
  wire  _GEN_86 = delay >= 8'h2 & _T_1 & _GEN_22; // @[div.scala 50:22 60:44]
  wire  S_tmp_19 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_86; // @[div.scala 50:22 58:46]
  wire  _GEN_83 = delay >= 8'h2 & _T_1 & _GEN_19; // @[div.scala 50:22 60:44]
  wire  S_tmp_16 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_83; // @[div.scala 50:22 58:46]
  wire  _GEN_84 = delay >= 8'h2 & _T_1 & _GEN_20; // @[div.scala 50:22 60:44]
  wire  S_tmp_17 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_84; // @[div.scala 50:22 58:46]
  wire [15:0] S_hi_lo = {S_tmp_16,S_tmp_17,S_tmp_18,S_tmp_19,S_tmp_20,S_tmp_21,S_tmp_22,S_tmp_23,S_hi_lo_lo}; // @[Cat.scala 31:58]
  wire  _GEN_81 = delay >= 8'h2 & _T_1 & _GEN_17; // @[div.scala 50:22 60:44]
  wire  S_tmp_14 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_81; // @[div.scala 50:22 58:46]
  wire  _GEN_82 = delay >= 8'h2 & _T_1 & _GEN_18; // @[div.scala 50:22 60:44]
  wire  S_tmp_15 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_82; // @[div.scala 50:22 58:46]
  wire  _GEN_79 = delay >= 8'h2 & _T_1 & _GEN_15; // @[div.scala 50:22 60:44]
  wire  S_tmp_12 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_79; // @[div.scala 50:22 58:46]
  wire  _GEN_80 = delay >= 8'h2 & _T_1 & _GEN_16; // @[div.scala 50:22 60:44]
  wire  S_tmp_13 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_80; // @[div.scala 50:22 58:46]
  wire  _GEN_77 = delay >= 8'h2 & _T_1 & _GEN_13; // @[div.scala 50:22 60:44]
  wire  S_tmp_10 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_77; // @[div.scala 50:22 58:46]
  wire  _GEN_78 = delay >= 8'h2 & _T_1 & _GEN_14; // @[div.scala 50:22 60:44]
  wire  S_tmp_11 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_78; // @[div.scala 50:22 58:46]
  wire  _GEN_75 = delay >= 8'h2 & _T_1 & _GEN_11; // @[div.scala 50:22 60:44]
  wire  S_tmp_8 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_75; // @[div.scala 50:22 58:46]
  wire  _GEN_76 = delay >= 8'h2 & _T_1 & _GEN_12; // @[div.scala 50:22 60:44]
  wire  S_tmp_9 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_76; // @[div.scala 50:22 58:46]
  wire [7:0] S_hi_hi_lo = {S_tmp_8,S_tmp_9,S_tmp_10,S_tmp_11,S_tmp_12,S_tmp_13,S_tmp_14,S_tmp_15}; // @[Cat.scala 31:58]
  wire  _GEN_73 = delay >= 8'h2 & _T_1 & _GEN_9; // @[div.scala 50:22 60:44]
  wire  S_tmp_6 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_73; // @[div.scala 50:22 58:46]
  wire  _GEN_74 = delay >= 8'h2 & _T_1 & _GEN_10; // @[div.scala 50:22 60:44]
  wire  S_tmp_7 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_74; // @[div.scala 50:22 58:46]
  wire  _GEN_71 = delay >= 8'h2 & _T_1 & _GEN_7; // @[div.scala 50:22 60:44]
  wire  S_tmp_4 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_71; // @[div.scala 50:22 58:46]
  wire  _GEN_72 = delay >= 8'h2 & _T_1 & _GEN_8; // @[div.scala 50:22 60:44]
  wire  S_tmp_5 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_72; // @[div.scala 50:22 58:46]
  wire  _GEN_69 = delay >= 8'h2 & _T_1 & _GEN_5; // @[div.scala 50:22 60:44]
  wire  S_tmp_2 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_69; // @[div.scala 50:22 58:46]
  wire  _GEN_70 = delay >= 8'h2 & _T_1 & _GEN_6; // @[div.scala 50:22 60:44]
  wire  S_tmp_3 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_70; // @[div.scala 50:22 58:46]
  wire  _GEN_67 = delay >= 8'h2 & _T_1 & _GEN_3; // @[div.scala 50:22 60:44]
  wire  S_tmp_0 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_67; // @[div.scala 50:22 58:46]
  wire  _GEN_68 = delay >= 8'h2 & _T_1 & _GEN_4; // @[div.scala 50:22 60:44]
  wire  S_tmp_1 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_68; // @[div.scala 50:22 58:46]
  wire [31:0] S_hi = {S_tmp_0,S_tmp_1,S_tmp_2,S_tmp_3,S_tmp_4,S_tmp_5,S_tmp_6,S_tmp_7,S_hi_hi_lo,S_hi_lo}; // @[Cat.scala 31:58]
  wire [63:0] _S_T = {S_hi,S_lo}; // @[Cat.scala 31:58]
  wire [63:0] _S_T_1 = _S_T | S; // @[div.scala 64:21]
  wire [128:0] _GEN_131 = delay >= 8'h2 & _T_1 ? _A_T_13 : {{1'd0}, _A_T}; // @[div.scala 60:44 54:5 62:7]
  wire [128:0] _GEN_199 = delay < 8'h2 & ~io_out_valid & start ? {{1'd0}, _A_T} : _GEN_131; // @[div.scala 58:46 54:5]
  wire  _GEN_202 = io_div_valid | start; // @[div.scala 66:21 67:11 23:25]
  wire [1:0] _clear_T_1 = clear + 2'h1; // @[div.scala 77:20]
  wire [128:0] _GEN_210 = clear == 2'h1 ? 129'h0 : _GEN_199; // @[div.scala 79:22 83:7]
  wire [63:0] _io_quotient_T_1 = ~S; // @[div.scala 92:47]
  wire [63:0] _io_quotient_T_3 = _io_quotient_T_1 + 64'h1; // @[div.scala 92:51]
  wire [63:0] _io_remainder_T_2 = ~A[127:64]; // @[div.scala 93:47]
  wire [63:0] _io_remainder_T_4 = _io_remainder_T_2 + 64'h1; // @[div.scala 93:64]
  wire [128:0] _GEN_280 = reset ? 129'h0 : _GEN_210; // @[div.scala 48:{18,18}]
  assign io_out_valid = cnt == 8'h40 & start; // @[div.scala 71:24]
  assign io_quotient = quotient_sign ? _io_quotient_T_3 : S; // @[div.scala 92:22]
  assign io_remainder = remainder_sign ? _io_remainder_T_4 : A[127:64]; // @[div.scala 93:22]
  always @(posedge clock) begin
    if (clear == 2'h1) begin // @[div.scala 79:22]
      dividend_reg <= 64'h0; // @[div.scala 86:18]
    end else if (start) begin // @[div.scala 33:14]
      if (io_div_signed & io_dividend[63]) begin // @[div.scala 31:18]
        dividend_reg <= _dividend_T_5;
      end else begin
        dividend_reg <= io_dividend;
      end
    end
    if (clear == 2'h1) begin // @[div.scala 79:22]
      divisor_reg <= 64'h0; // @[div.scala 87:18]
    end else if (start) begin // @[div.scala 33:14]
      if (io_div_signed & io_divisor[63]) begin // @[div.scala 32:18]
        divisor_reg <= _divisor_T_5;
      end else begin
        divisor_reg <= io_divisor;
      end
    end
    if (reset) begin // @[div.scala 23:25]
      start <= 1'h0; // @[div.scala 23:25]
    end else if (cnt == 8'h40 & start) begin // @[div.scala 71:33]
      start <= 1'h0; // @[div.scala 72:11]
    end else begin
      start <= _GEN_202;
    end
    if (reset) begin // @[div.scala 25:24]
      delay <= 8'h0; // @[div.scala 25:24]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      delay <= 8'h0; // @[div.scala 88:11]
    end else if (delay < 8'h2 & ~io_out_valid & start) begin // @[div.scala 58:46]
      delay <= _delay_T_1; // @[div.scala 59:11]
    end
    if (reset) begin // @[div.scala 27:24]
      clear <= 2'h0; // @[div.scala 27:24]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      clear <= 2'h0; // @[div.scala 89:11]
    end else if (io_out_valid) begin // @[div.scala 76:21]
      clear <= _clear_T_1; // @[div.scala 77:11]
    end
    if (reset) begin // @[div.scala 42:31]
      quotient_sign <= 1'h0; // @[div.scala 42:31]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      quotient_sign <= 1'h0; // @[div.scala 81:20]
    end else if (io_div_valid) begin // @[div.scala 44:24]
      quotient_sign <= io_div_signed & (io_dividend[63] ^ io_divisor[63]);
    end else begin
      quotient_sign <= remainder_sign;
    end
    if (reset) begin // @[div.scala 43:31]
      remainder_sign <= 1'h0; // @[div.scala 43:31]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      remainder_sign <= 1'h0; // @[div.scala 82:20]
    end else if (io_div_valid) begin // @[div.scala 45:24]
      remainder_sign <= _dividend_T_1;
    end
    A <= _GEN_280[127:0]; // @[div.scala 48:{18,18}]
    if (reset) begin // @[div.scala 49:18]
      B <= 64'h0; // @[div.scala 49:18]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      B <= 64'h0; // @[div.scala 84:7]
    end else begin
      B <= divisor_reg; // @[div.scala 55:5]
    end
    if (reset) begin // @[div.scala 51:18]
      S <= 64'h0; // @[div.scala 51:18]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      S <= 64'h0; // @[div.scala 85:7]
    end else if (!(delay < 8'h2 & ~io_out_valid & start)) begin // @[div.scala 58:46]
      if (delay >= 8'h2 & _T_1) begin // @[div.scala 60:44]
        S <= _S_T_1; // @[div.scala 64:7]
      end
    end
    if (reset) begin // @[div.scala 52:20]
      cnt <= 8'h0; // @[div.scala 52:20]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      cnt <= 8'h0; // @[div.scala 80:9]
    end else if (!(delay < 8'h2 & ~io_out_valid & start)) begin // @[div.scala 58:46]
      if (delay >= 8'h2 & _T_1) begin // @[div.scala 60:44]
        cnt <= _cnt_T_1; // @[div.scala 63:9]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  dividend_reg = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  divisor_reg = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  start = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  delay = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  clear = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  quotient_sign = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  remainder_sign = _RAND_6[0:0];
  _RAND_7 = {4{`RANDOM}};
  A = _RAND_7[127:0];
  _RAND_8 = {2{`RANDOM}};
  B = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  S = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  cnt = _RAND_10[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module div_1(
  input         clock,
  input         reset,
  input  [31:0] io_dividend,
  input  [31:0] io_divisor,
  input         io_div_valid,
  input         io_div_signed,
  output        io_out_valid,
  output [31:0] io_quotient,
  output [31:0] io_remainder
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] dividend_reg; // @[div.scala 21:25]
  reg [31:0] divisor_reg; // @[div.scala 22:25]
  reg  start; // @[div.scala 23:25]
  reg [7:0] delay; // @[div.scala 25:24]
  reg [1:0] clear; // @[div.scala 27:24]
  wire  _dividend_T_1 = io_div_signed & io_dividend[31]; // @[div.scala 31:34]
  wire [31:0] _dividend_T_3 = ~io_dividend; // @[div.scala 31:66]
  wire [31:0] _dividend_T_5 = _dividend_T_3 + 32'h1; // @[div.scala 31:80]
  wire [31:0] _divisor_T_3 = ~io_divisor; // @[div.scala 32:65]
  wire [31:0] _divisor_T_5 = _divisor_T_3 + 32'h1; // @[div.scala 32:78]
  reg  quotient_sign; // @[div.scala 42:31]
  reg  remainder_sign; // @[div.scala 43:31]
  reg [63:0] A; // @[div.scala 48:18]
  reg [31:0] B; // @[div.scala 49:18]
  reg [31:0] S; // @[div.scala 51:18]
  reg [7:0] cnt; // @[div.scala 52:20]
  wire [63:0] _A_T = {32'h0,dividend_reg}; // @[Cat.scala 31:58]
  wire  _T_1 = ~io_out_valid; // @[div.scala 58:23]
  wire [7:0] _delay_T_1 = delay + 8'h1; // @[div.scala 59:20]
  wire [32:0] _S_tmp_T_1 = {1'h0,B}; // @[Cat.scala 31:58]
  wire  _S_tmp_T_2 = A[63:31] >= _S_tmp_T_1; // @[div.scala 61:42]
  wire  _GEN_3 = 5'h0 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_4 = 5'h1 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_5 = 5'h2 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_6 = 5'h3 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_7 = 5'h4 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_8 = 5'h5 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_9 = 5'h6 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_10 = 5'h7 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_11 = 5'h8 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_12 = 5'h9 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_13 = 5'ha == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_14 = 5'hb == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_15 = 5'hc == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_16 = 5'hd == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_17 = 5'he == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_18 = 5'hf == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_19 = 5'h10 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_20 = 5'h11 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_21 = 5'h12 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_22 = 5'h13 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_23 = 5'h14 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_24 = 5'h15 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_25 = 5'h16 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_26 = 5'h17 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_27 = 5'h18 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_28 = 5'h19 == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_29 = 5'h1a == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_30 = 5'h1b == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_31 = 5'h1c == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_32 = 5'h1d == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_33 = 5'h1e == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire  _GEN_34 = 5'h1f == cnt[4:0] & A[63:31] >= _S_tmp_T_1; // @[div.scala 61:{16,16} 50:22]
  wire [63:0] _A_T_5 = {33'h0,A[30:0]}; // @[Cat.scala 31:58]
  wire [32:0] _A_T_9 = A[63:31] - _S_tmp_T_1; // @[div.scala 62:106]
  wire [63:0] _A_T_10 = {_A_T_9, 31'h0}; // @[div.scala 62:121]
  wire [63:0] _A_T_11 = _A_T_5 | _A_T_10; // @[div.scala 62:84]
  wire [63:0] _A_T_12 = _S_tmp_T_2 ? _A_T_11 : A; // @[div.scala 62:14]
  wire [64:0] _A_T_13 = {_A_T_12, 1'h0}; // @[div.scala 62:137]
  wire [7:0] _cnt_T_1 = cnt + 8'h1; // @[div.scala 63:16]
  wire  _GEN_65 = delay >= 8'h2 & _T_1 & _GEN_33; // @[div.scala 50:22 60:44]
  wire  S_tmp_30 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_65; // @[div.scala 50:22 58:46]
  wire  _GEN_66 = delay >= 8'h2 & _T_1 & _GEN_34; // @[div.scala 50:22 60:44]
  wire  S_tmp_31 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_66; // @[div.scala 50:22 58:46]
  wire  _GEN_63 = delay >= 8'h2 & _T_1 & _GEN_31; // @[div.scala 50:22 60:44]
  wire  S_tmp_28 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_63; // @[div.scala 50:22 58:46]
  wire  _GEN_64 = delay >= 8'h2 & _T_1 & _GEN_32; // @[div.scala 50:22 60:44]
  wire  S_tmp_29 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_64; // @[div.scala 50:22 58:46]
  wire  _GEN_61 = delay >= 8'h2 & _T_1 & _GEN_29; // @[div.scala 50:22 60:44]
  wire  S_tmp_26 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_61; // @[div.scala 50:22 58:46]
  wire  _GEN_62 = delay >= 8'h2 & _T_1 & _GEN_30; // @[div.scala 50:22 60:44]
  wire  S_tmp_27 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_62; // @[div.scala 50:22 58:46]
  wire  _GEN_59 = delay >= 8'h2 & _T_1 & _GEN_27; // @[div.scala 50:22 60:44]
  wire  S_tmp_24 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_59; // @[div.scala 50:22 58:46]
  wire  _GEN_60 = delay >= 8'h2 & _T_1 & _GEN_28; // @[div.scala 50:22 60:44]
  wire  S_tmp_25 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_60; // @[div.scala 50:22 58:46]
  wire [7:0] S_lo_lo = {S_tmp_24,S_tmp_25,S_tmp_26,S_tmp_27,S_tmp_28,S_tmp_29,S_tmp_30,S_tmp_31}; // @[Cat.scala 31:58]
  wire  _GEN_57 = delay >= 8'h2 & _T_1 & _GEN_25; // @[div.scala 50:22 60:44]
  wire  S_tmp_22 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_57; // @[div.scala 50:22 58:46]
  wire  _GEN_58 = delay >= 8'h2 & _T_1 & _GEN_26; // @[div.scala 50:22 60:44]
  wire  S_tmp_23 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_58; // @[div.scala 50:22 58:46]
  wire  _GEN_55 = delay >= 8'h2 & _T_1 & _GEN_23; // @[div.scala 50:22 60:44]
  wire  S_tmp_20 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_55; // @[div.scala 50:22 58:46]
  wire  _GEN_56 = delay >= 8'h2 & _T_1 & _GEN_24; // @[div.scala 50:22 60:44]
  wire  S_tmp_21 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_56; // @[div.scala 50:22 58:46]
  wire  _GEN_53 = delay >= 8'h2 & _T_1 & _GEN_21; // @[div.scala 50:22 60:44]
  wire  S_tmp_18 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_53; // @[div.scala 50:22 58:46]
  wire  _GEN_54 = delay >= 8'h2 & _T_1 & _GEN_22; // @[div.scala 50:22 60:44]
  wire  S_tmp_19 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_54; // @[div.scala 50:22 58:46]
  wire  _GEN_51 = delay >= 8'h2 & _T_1 & _GEN_19; // @[div.scala 50:22 60:44]
  wire  S_tmp_16 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_51; // @[div.scala 50:22 58:46]
  wire  _GEN_52 = delay >= 8'h2 & _T_1 & _GEN_20; // @[div.scala 50:22 60:44]
  wire  S_tmp_17 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_52; // @[div.scala 50:22 58:46]
  wire [15:0] S_lo = {S_tmp_16,S_tmp_17,S_tmp_18,S_tmp_19,S_tmp_20,S_tmp_21,S_tmp_22,S_tmp_23,S_lo_lo}; // @[Cat.scala 31:58]
  wire  _GEN_49 = delay >= 8'h2 & _T_1 & _GEN_17; // @[div.scala 50:22 60:44]
  wire  S_tmp_14 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_49; // @[div.scala 50:22 58:46]
  wire  _GEN_50 = delay >= 8'h2 & _T_1 & _GEN_18; // @[div.scala 50:22 60:44]
  wire  S_tmp_15 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_50; // @[div.scala 50:22 58:46]
  wire  _GEN_47 = delay >= 8'h2 & _T_1 & _GEN_15; // @[div.scala 50:22 60:44]
  wire  S_tmp_12 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_47; // @[div.scala 50:22 58:46]
  wire  _GEN_48 = delay >= 8'h2 & _T_1 & _GEN_16; // @[div.scala 50:22 60:44]
  wire  S_tmp_13 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_48; // @[div.scala 50:22 58:46]
  wire  _GEN_45 = delay >= 8'h2 & _T_1 & _GEN_13; // @[div.scala 50:22 60:44]
  wire  S_tmp_10 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_45; // @[div.scala 50:22 58:46]
  wire  _GEN_46 = delay >= 8'h2 & _T_1 & _GEN_14; // @[div.scala 50:22 60:44]
  wire  S_tmp_11 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_46; // @[div.scala 50:22 58:46]
  wire  _GEN_43 = delay >= 8'h2 & _T_1 & _GEN_11; // @[div.scala 50:22 60:44]
  wire  S_tmp_8 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_43; // @[div.scala 50:22 58:46]
  wire  _GEN_44 = delay >= 8'h2 & _T_1 & _GEN_12; // @[div.scala 50:22 60:44]
  wire  S_tmp_9 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_44; // @[div.scala 50:22 58:46]
  wire [7:0] S_hi_lo = {S_tmp_8,S_tmp_9,S_tmp_10,S_tmp_11,S_tmp_12,S_tmp_13,S_tmp_14,S_tmp_15}; // @[Cat.scala 31:58]
  wire  _GEN_41 = delay >= 8'h2 & _T_1 & _GEN_9; // @[div.scala 50:22 60:44]
  wire  S_tmp_6 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_41; // @[div.scala 50:22 58:46]
  wire  _GEN_42 = delay >= 8'h2 & _T_1 & _GEN_10; // @[div.scala 50:22 60:44]
  wire  S_tmp_7 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_42; // @[div.scala 50:22 58:46]
  wire  _GEN_39 = delay >= 8'h2 & _T_1 & _GEN_7; // @[div.scala 50:22 60:44]
  wire  S_tmp_4 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_39; // @[div.scala 50:22 58:46]
  wire  _GEN_40 = delay >= 8'h2 & _T_1 & _GEN_8; // @[div.scala 50:22 60:44]
  wire  S_tmp_5 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_40; // @[div.scala 50:22 58:46]
  wire  _GEN_37 = delay >= 8'h2 & _T_1 & _GEN_5; // @[div.scala 50:22 60:44]
  wire  S_tmp_2 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_37; // @[div.scala 50:22 58:46]
  wire  _GEN_38 = delay >= 8'h2 & _T_1 & _GEN_6; // @[div.scala 50:22 60:44]
  wire  S_tmp_3 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_38; // @[div.scala 50:22 58:46]
  wire  _GEN_35 = delay >= 8'h2 & _T_1 & _GEN_3; // @[div.scala 50:22 60:44]
  wire  S_tmp_0 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_35; // @[div.scala 50:22 58:46]
  wire  _GEN_36 = delay >= 8'h2 & _T_1 & _GEN_4; // @[div.scala 50:22 60:44]
  wire  S_tmp_1 = delay < 8'h2 & ~io_out_valid & start ? 1'h0 : _GEN_36; // @[div.scala 50:22 58:46]
  wire [31:0] _S_T = {S_tmp_0,S_tmp_1,S_tmp_2,S_tmp_3,S_tmp_4,S_tmp_5,S_tmp_6,S_tmp_7,S_hi_lo,S_lo}; // @[Cat.scala 31:58]
  wire [31:0] _S_T_1 = _S_T | S; // @[div.scala 64:21]
  wire [64:0] _GEN_67 = delay >= 8'h2 & _T_1 ? _A_T_13 : {{1'd0}, _A_T}; // @[div.scala 60:44 54:5 62:7]
  wire [64:0] _GEN_103 = delay < 8'h2 & ~io_out_valid & start ? {{1'd0}, _A_T} : _GEN_67; // @[div.scala 58:46 54:5]
  wire  _GEN_106 = io_div_valid | start; // @[div.scala 66:21 67:11 23:25]
  wire [1:0] _clear_T_1 = clear + 2'h1; // @[div.scala 77:20]
  wire [64:0] _GEN_114 = clear == 2'h1 ? 65'h0 : _GEN_103; // @[div.scala 79:22 83:7]
  wire [31:0] _io_quotient_T_1 = ~S; // @[div.scala 92:47]
  wire [31:0] _io_quotient_T_3 = _io_quotient_T_1 + 32'h1; // @[div.scala 92:51]
  wire [31:0] _io_remainder_T_2 = ~A[63:32]; // @[div.scala 93:47]
  wire [31:0] _io_remainder_T_4 = _io_remainder_T_2 + 32'h1; // @[div.scala 93:64]
  wire [64:0] _GEN_152 = reset ? 65'h0 : _GEN_114; // @[div.scala 48:{18,18}]
  assign io_out_valid = cnt == 8'h20 & start; // @[div.scala 71:24]
  assign io_quotient = quotient_sign ? _io_quotient_T_3 : S; // @[div.scala 92:22]
  assign io_remainder = remainder_sign ? _io_remainder_T_4 : A[63:32]; // @[div.scala 93:22]
  always @(posedge clock) begin
    if (clear == 2'h1) begin // @[div.scala 79:22]
      dividend_reg <= 32'h0; // @[div.scala 86:18]
    end else if (start) begin // @[div.scala 33:14]
      if (io_div_signed & io_dividend[31]) begin // @[div.scala 31:18]
        dividend_reg <= _dividend_T_5;
      end else begin
        dividend_reg <= io_dividend;
      end
    end
    if (clear == 2'h1) begin // @[div.scala 79:22]
      divisor_reg <= 32'h0; // @[div.scala 87:18]
    end else if (start) begin // @[div.scala 33:14]
      if (io_div_signed & io_divisor[31]) begin // @[div.scala 32:18]
        divisor_reg <= _divisor_T_5;
      end else begin
        divisor_reg <= io_divisor;
      end
    end
    if (reset) begin // @[div.scala 23:25]
      start <= 1'h0; // @[div.scala 23:25]
    end else if (cnt == 8'h20 & start) begin // @[div.scala 71:33]
      start <= 1'h0; // @[div.scala 72:11]
    end else begin
      start <= _GEN_106;
    end
    if (reset) begin // @[div.scala 25:24]
      delay <= 8'h0; // @[div.scala 25:24]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      delay <= 8'h0; // @[div.scala 88:11]
    end else if (delay < 8'h2 & ~io_out_valid & start) begin // @[div.scala 58:46]
      delay <= _delay_T_1; // @[div.scala 59:11]
    end
    if (reset) begin // @[div.scala 27:24]
      clear <= 2'h0; // @[div.scala 27:24]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      clear <= 2'h0; // @[div.scala 89:11]
    end else if (io_out_valid) begin // @[div.scala 76:21]
      clear <= _clear_T_1; // @[div.scala 77:11]
    end
    if (reset) begin // @[div.scala 42:31]
      quotient_sign <= 1'h0; // @[div.scala 42:31]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      quotient_sign <= 1'h0; // @[div.scala 81:20]
    end else if (io_div_valid) begin // @[div.scala 44:24]
      quotient_sign <= io_div_signed & (io_dividend[31] ^ io_divisor[31]);
    end else begin
      quotient_sign <= remainder_sign;
    end
    if (reset) begin // @[div.scala 43:31]
      remainder_sign <= 1'h0; // @[div.scala 43:31]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      remainder_sign <= 1'h0; // @[div.scala 82:20]
    end else if (io_div_valid) begin // @[div.scala 45:24]
      remainder_sign <= _dividend_T_1;
    end
    A <= _GEN_152[63:0]; // @[div.scala 48:{18,18}]
    if (reset) begin // @[div.scala 49:18]
      B <= 32'h0; // @[div.scala 49:18]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      B <= 32'h0; // @[div.scala 84:7]
    end else begin
      B <= divisor_reg; // @[div.scala 55:5]
    end
    if (reset) begin // @[div.scala 51:18]
      S <= 32'h0; // @[div.scala 51:18]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      S <= 32'h0; // @[div.scala 85:7]
    end else if (!(delay < 8'h2 & ~io_out_valid & start)) begin // @[div.scala 58:46]
      if (delay >= 8'h2 & _T_1) begin // @[div.scala 60:44]
        S <= _S_T_1; // @[div.scala 64:7]
      end
    end
    if (reset) begin // @[div.scala 52:20]
      cnt <= 8'h0; // @[div.scala 52:20]
    end else if (clear == 2'h1) begin // @[div.scala 79:22]
      cnt <= 8'h0; // @[div.scala 80:9]
    end else if (!(delay < 8'h2 & ~io_out_valid & start)) begin // @[div.scala 58:46]
      if (delay >= 8'h2 & _T_1) begin // @[div.scala 60:44]
        cnt <= _cnt_T_1; // @[div.scala 63:9]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dividend_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  divisor_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  start = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  delay = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  clear = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  quotient_sign = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  remainder_sign = _RAND_6[0:0];
  _RAND_7 = {2{`RANDOM}};
  A = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  B = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  S = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  cnt = _RAND_10[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EXU(
  input         clock,
  input         reset,
  input         io_ms_allowin,
  output        io_es_allowin,
  input         io_ds_to_es_valid,
  output        io_es_to_ms_valid,
  input  [7:0]  io_de_bus_OP,
  input         io_de_bus_res_from_mem,
  input         io_de_bus_gr_we,
  input         io_de_bus_MemWen,
  input  [7:0]  io_de_bus_wmask,
  input  [31:0] io_de_bus_ds_pc,
  input  [4:0]  io_de_bus_dest,
  input  [63:0] io_de_bus_imm,
  input  [63:0] io_de_bus_rdata1,
  input  [63:0] io_de_bus_rdata2,
  input  [2:0]  io_de_bus_ld_type,
  input  [31:0] io_de_bus_inst,
  input  [63:0] io_de_bus_csr_rdata,
  input  [2:0]  io_de_bus_csr_waddr1,
  input  [2:0]  io_de_bus_csr_waddr2,
  input         io_de_bus_csr_wen,
  input         io_de_bus_eval,
  input         io_de_bus_is_ld,
  output        io_em_bus_res_from_mem,
  output        io_em_bus_gr_we,
  output [4:0]  io_em_bus_dest,
  output [63:0] io_em_bus_alu_result,
  output [31:0] io_em_bus_ex_pc,
  output [2:0]  io_em_bus_ld_type,
  output [31:0] io_em_bus_inst,
  output [63:0] io_em_bus_csr_wdata,
  output        io_em_bus_csr_wen,
  output [2:0]  io_em_bus_csr_waddr1,
  output [2:0]  io_em_bus_csr_waddr2,
  output        io_em_bus_eval,
  output        io_em_bus_is_ld,
  output        io_em_bus_MemWen,
  output [63:0] io_em_bus_Memwdata,
  output [7:0]  io_em_bus_wmask,
  output        io_es_dest_valid_gr_we,
  output        io_es_dest_valid_es_valid,
  output [4:0]  io_es_dest_valid_dest,
  output [63:0] io_es_dest_valid_es_forward_data,
  output        io_es_dest_valid_es_is_ld,
  output        io_es_dest_valid_es_ready_go,
  output        io_es_dest_valid_es_to_ms_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire  mul_clock; // @[EXU.scala 51:23]
  wire  mul_reset; // @[EXU.scala 51:23]
  wire  mul_io_mul_valid; // @[EXU.scala 51:23]
  wire [63:0] mul_io_multiplicand; // @[EXU.scala 51:23]
  wire [63:0] mul_io_multiplier; // @[EXU.scala 51:23]
  wire  mul_io_out_valid; // @[EXU.scala 51:23]
  wire [63:0] mul_io_result_lo; // @[EXU.scala 51:23]
  wire  mul_1_clock; // @[EXU.scala 52:23]
  wire  mul_1_reset; // @[EXU.scala 52:23]
  wire  mul_1_io_mul_valid; // @[EXU.scala 52:23]
  wire [31:0] mul_1_io_multiplicand; // @[EXU.scala 52:23]
  wire [31:0] mul_1_io_multiplier; // @[EXU.scala 52:23]
  wire  mul_1_io_out_valid; // @[EXU.scala 52:23]
  wire [31:0] mul_1_io_result_lo; // @[EXU.scala 52:23]
  wire  div_clock; // @[EXU.scala 70:23]
  wire  div_reset; // @[EXU.scala 70:23]
  wire [63:0] div_io_dividend; // @[EXU.scala 70:23]
  wire [63:0] div_io_divisor; // @[EXU.scala 70:23]
  wire  div_io_div_valid; // @[EXU.scala 70:23]
  wire  div_io_div_signed; // @[EXU.scala 70:23]
  wire  div_io_out_valid; // @[EXU.scala 70:23]
  wire [63:0] div_io_quotient; // @[EXU.scala 70:23]
  wire [63:0] div_io_remainder; // @[EXU.scala 70:23]
  wire  div_1_clock; // @[EXU.scala 71:23]
  wire  div_1_reset; // @[EXU.scala 71:23]
  wire [31:0] div_1_io_dividend; // @[EXU.scala 71:23]
  wire [31:0] div_1_io_divisor; // @[EXU.scala 71:23]
  wire  div_1_io_div_valid; // @[EXU.scala 71:23]
  wire  div_1_io_div_signed; // @[EXU.scala 71:23]
  wire  div_1_io_out_valid; // @[EXU.scala 71:23]
  wire [31:0] div_1_io_quotient; // @[EXU.scala 71:23]
  wire [31:0] div_1_io_remainder; // @[EXU.scala 71:23]
  reg [7:0] de_bus_r_OP; // @[EXU.scala 23:28]
  reg  de_bus_r_res_from_mem; // @[EXU.scala 23:28]
  reg  de_bus_r_gr_we; // @[EXU.scala 23:28]
  reg  de_bus_r_MemWen; // @[EXU.scala 23:28]
  reg [7:0] de_bus_r_wmask; // @[EXU.scala 23:28]
  reg [31:0] de_bus_r_ds_pc; // @[EXU.scala 23:28]
  reg [4:0] de_bus_r_dest; // @[EXU.scala 23:28]
  reg [63:0] de_bus_r_imm; // @[EXU.scala 23:28]
  reg [63:0] de_bus_r_rdata1; // @[EXU.scala 23:28]
  reg [63:0] de_bus_r_rdata2; // @[EXU.scala 23:28]
  reg [2:0] de_bus_r_ld_type; // @[EXU.scala 23:28]
  reg [31:0] de_bus_r_inst; // @[EXU.scala 23:28]
  reg [63:0] de_bus_r_csr_rdata; // @[EXU.scala 23:28]
  reg [2:0] de_bus_r_csr_waddr1; // @[EXU.scala 23:28]
  reg [2:0] de_bus_r_csr_waddr2; // @[EXU.scala 23:28]
  reg  de_bus_r_csr_wen; // @[EXU.scala 23:28]
  reg  de_bus_r_eval; // @[EXU.scala 23:28]
  reg  de_bus_r_is_ld; // @[EXU.scala 23:28]
  reg  es_valid; // @[EXU.scala 24:28]
  wire  is_mul_64 = de_bus_r_OP == 8'h4; // @[EXU.scala 53:31]
  wire  is_mul_32 = de_bus_r_OP == 8'h5; // @[EXU.scala 54:31]
  wire  _is_div_64_T = de_bus_r_OP == 8'h6; // @[EXU.scala 72:32]
  wire  is_div_64 = de_bus_r_OP == 8'h6 | de_bus_r_OP == 8'h7; // @[EXU.scala 72:44]
  wire  _is_div_32_T = de_bus_r_OP == 8'h8; // @[EXU.scala 73:32]
  wire  is_div_32 = de_bus_r_OP == 8'h8 | de_bus_r_OP == 8'h9; // @[EXU.scala 73:45]
  wire  _is_rem_64_T = de_bus_r_OP == 8'h15; // @[EXU.scala 74:32]
  wire  is_rem_64 = de_bus_r_OP == 8'h15 | de_bus_r_OP == 8'h16; // @[EXU.scala 74:44]
  wire  _is_rem_32_T = de_bus_r_OP == 8'h17; // @[EXU.scala 75:32]
  wire  is_rem_32 = de_bus_r_OP == 8'h17 | de_bus_r_OP == 8'h18; // @[EXU.scala 75:45]
  wire [63:0] _result_T_1 = de_bus_r_rdata1 + de_bus_r_rdata2; // @[EXU.scala 96:24]
  wire [31:0] _result_T_5 = de_bus_r_rdata1[31:0] + de_bus_r_rdata2[31:0]; // @[EXU.scala 97:37]
  wire [31:0] _result_T_8 = _result_T_5[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _result_T_10 = {_result_T_8,_result_T_5}; // @[Cat.scala 31:58]
  wire [63:0] _result_T_12 = de_bus_r_rdata1 - de_bus_r_rdata2; // @[EXU.scala 98:24]
  wire [31:0] _result_T_16 = de_bus_r_rdata1[31:0] - de_bus_r_rdata2[31:0]; // @[EXU.scala 99:36]
  wire [31:0] _result_T_19 = _result_T_16[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _result_T_21 = {_result_T_19,_result_T_16}; // @[Cat.scala 31:58]
  wire [31:0] _result_T_24 = mul_1_io_result_lo[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _result_T_25 = mul_1_io_result_lo; // @[EXU.scala 43:66]
  wire [63:0] _result_T_26 = {_result_T_24,_result_T_25}; // @[Cat.scala 31:58]
  wire [31:0] _result_T_29 = div_1_io_quotient[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _result_T_30 = div_1_io_quotient; // @[EXU.scala 43:66]
  wire [63:0] _result_T_31 = {_result_T_29,_result_T_30}; // @[Cat.scala 31:58]
  wire [126:0] _GEN_7 = {{63'd0}, de_bus_r_rdata1}; // @[EXU.scala 106:24]
  wire [126:0] _result_T_38 = _GEN_7 << de_bus_r_rdata2[5:0]; // @[EXU.scala 106:24]
  wire  _result_T_41 = $signed(de_bus_r_rdata1) < $signed(de_bus_r_rdata2); // @[EXU.scala 107:35]
  wire  _result_T_43 = de_bus_r_rdata1 < de_bus_r_rdata2; // @[EXU.scala 108:29]
  wire [62:0] _GEN_15 = {{31'd0}, de_bus_r_rdata1[31:0]}; // @[EXU.scala 109:37]
  wire [62:0] _result_T_47 = _GEN_15 << de_bus_r_rdata2[4:0]; // @[EXU.scala 109:37]
  wire [31:0] _result_T_50 = _result_T_47[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _result_T_52 = {_result_T_50,_result_T_47[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _result_T_56 = $signed(de_bus_r_rdata1) >>> de_bus_r_rdata2[5:0]; // @[EXU.scala 110:46]
  wire [31:0] _result_T_58 = de_bus_r_rdata1[31:0]; // @[EXU.scala 111:37]
  wire [31:0] _result_T_61 = $signed(_result_T_58) >>> de_bus_r_rdata2[4:0]; // @[EXU.scala 111:59]
  wire [31:0] _result_T_64 = _result_T_61[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _result_T_66 = {_result_T_64,_result_T_61}; // @[Cat.scala 31:58]
  wire [63:0] _result_T_68 = de_bus_r_rdata1 >> de_bus_r_rdata2[5:0]; // @[EXU.scala 112:24]
  wire [31:0] _result_T_71 = de_bus_r_rdata1[31:0] >> de_bus_r_rdata2[4:0]; // @[EXU.scala 113:37]
  wire [31:0] _result_T_74 = _result_T_71[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _result_T_76 = {_result_T_74,_result_T_71}; // @[Cat.scala 31:58]
  wire [63:0] _result_T_77 = de_bus_r_rdata1 ^ de_bus_r_rdata2; // @[EXU.scala 114:24]
  wire [63:0] _result_T_78 = de_bus_r_rdata1 & de_bus_r_rdata2; // @[EXU.scala 115:24]
  wire [63:0] _result_T_79 = de_bus_r_rdata1 | de_bus_r_rdata2; // @[EXU.scala 116:23]
  wire [31:0] _result_T_82 = div_1_io_remainder[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [31:0] _result_T_83 = div_1_io_remainder; // @[EXU.scala 43:66]
  wire [63:0] _result_T_84 = {_result_T_82,_result_T_83}; // @[Cat.scala 31:58]
  wire [63:0] _result_T_91 = de_bus_r_rdata1 + de_bus_r_imm; // @[EXU.scala 122:25]
  wire [63:0] _GEN_5 = {{32'd0}, de_bus_r_rdata1[31:0]}; // @[EXU.scala 123:38]
  wire [63:0] _result_T_94 = _GEN_5 + de_bus_r_imm; // @[EXU.scala 123:38]
  wire [31:0] _result_T_97 = _result_T_94[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _result_T_99 = {_result_T_97,_result_T_94[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] ex_pc = {{32'd0}, de_bus_r_ds_pc};
  wire [63:0] _result_T_101 = ex_pc + 64'h4; // @[EXU.scala 124:26]
  wire [126:0] _GEN_16 = {{63'd0}, de_bus_r_rdata1}; // @[EXU.scala 132:25]
  wire [126:0] _result_T_117 = _GEN_16 << de_bus_r_imm[5:0]; // @[EXU.scala 132:25]
  wire [62:0] _GEN_17 = {{31'd0}, de_bus_r_rdata1[31:0]}; // @[EXU.scala 133:39]
  wire [62:0] _result_T_120 = _GEN_17 << de_bus_r_imm[4:0]; // @[EXU.scala 133:39]
  wire [31:0] _result_T_123 = _result_T_120[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _result_T_125 = {_result_T_123,_result_T_120[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _result_T_127 = de_bus_r_rdata1 >> de_bus_r_imm[5:0]; // @[EXU.scala 134:25]
  wire [31:0] _result_T_130 = de_bus_r_rdata1[31:0] >> de_bus_r_imm[4:0]; // @[EXU.scala 135:39]
  wire [31:0] _result_T_133 = _result_T_130[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _result_T_135 = {_result_T_133,_result_T_130}; // @[Cat.scala 31:58]
  wire  _result_T_138 = $signed(de_bus_r_rdata1) < $signed(de_bus_r_imm); // @[EXU.scala 136:36]
  wire  _result_T_140 = de_bus_r_rdata1 < de_bus_r_imm; // @[EXU.scala 137:30]
  wire [63:0] _result_T_142 = de_bus_r_rdata1 & de_bus_r_imm; // @[EXU.scala 138:25]
  wire [63:0] _result_T_143 = de_bus_r_rdata1 ^ de_bus_r_imm; // @[EXU.scala 139:25]
  wire [63:0] _result_T_144 = de_bus_r_rdata1 | de_bus_r_imm; // @[EXU.scala 140:24]
  wire [63:0] _result_T_148 = $signed(de_bus_r_rdata1) >>> de_bus_r_imm[5:0]; // @[EXU.scala 141:46]
  wire [31:0] _result_T_153 = $signed(_result_T_58) >>> de_bus_r_imm[4:0]; // @[EXU.scala 142:60]
  wire [31:0] _result_T_156 = _result_T_153[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _result_T_158 = {_result_T_156,_result_T_153}; // @[Cat.scala 31:58]
  wire [63:0] _result_T_168 = ex_pc + de_bus_r_imm; // @[EXU.scala 153:27]
  wire [63:0] _result_T_172 = 8'h0 == de_bus_r_OP ? _result_T_1 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _result_T_174 = 8'h1 == de_bus_r_OP ? _result_T_10 : _result_T_172; // @[Mux.scala 81:58]
  wire [63:0] _result_T_176 = 8'h2 == de_bus_r_OP ? _result_T_12 : _result_T_174; // @[Mux.scala 81:58]
  wire [63:0] _result_T_178 = 8'h3 == de_bus_r_OP ? _result_T_21 : _result_T_176; // @[Mux.scala 81:58]
  wire [63:0] _result_T_180 = 8'h4 == de_bus_r_OP ? mul_io_result_lo : _result_T_178; // @[Mux.scala 81:58]
  wire [63:0] _result_T_182 = 8'h5 == de_bus_r_OP ? _result_T_26 : _result_T_180; // @[Mux.scala 81:58]
  wire [63:0] _result_T_184 = 8'h6 == de_bus_r_OP ? div_io_quotient : _result_T_182; // @[Mux.scala 81:58]
  wire [63:0] _result_T_186 = 8'h7 == de_bus_r_OP ? div_io_quotient : _result_T_184; // @[Mux.scala 81:58]
  wire [63:0] _result_T_188 = 8'h8 == de_bus_r_OP ? _result_T_31 : _result_T_186; // @[Mux.scala 81:58]
  wire [63:0] _result_T_190 = 8'h9 == de_bus_r_OP ? _result_T_31 : _result_T_188; // @[Mux.scala 81:58]
  wire [126:0] _result_T_192 = 8'ha == de_bus_r_OP ? _result_T_38 : {{63'd0}, _result_T_190}; // @[Mux.scala 81:58]
  wire [126:0] _result_T_194 = 8'hb == de_bus_r_OP ? {{126'd0}, _result_T_41} : _result_T_192; // @[Mux.scala 81:58]
  wire [126:0] _result_T_196 = 8'hc == de_bus_r_OP ? {{126'd0}, _result_T_43} : _result_T_194; // @[Mux.scala 81:58]
  wire [126:0] _result_T_198 = 8'hd == de_bus_r_OP ? {{63'd0}, _result_T_52} : _result_T_196; // @[Mux.scala 81:58]
  wire [126:0] _result_T_200 = 8'h13 == de_bus_r_OP ? {{63'd0}, _result_T_56} : _result_T_198; // @[Mux.scala 81:58]
  wire [126:0] _result_T_202 = 8'he == de_bus_r_OP ? {{63'd0}, _result_T_66} : _result_T_200; // @[Mux.scala 81:58]
  wire [126:0] _result_T_204 = 8'hf == de_bus_r_OP ? {{63'd0}, _result_T_68} : _result_T_202; // @[Mux.scala 81:58]
  wire [126:0] _result_T_206 = 8'h10 == de_bus_r_OP ? {{63'd0}, _result_T_76} : _result_T_204; // @[Mux.scala 81:58]
  wire [126:0] _result_T_208 = 8'h11 == de_bus_r_OP ? {{63'd0}, _result_T_77} : _result_T_206; // @[Mux.scala 81:58]
  wire [126:0] _result_T_210 = 8'h12 == de_bus_r_OP ? {{63'd0}, _result_T_78} : _result_T_208; // @[Mux.scala 81:58]
  wire [126:0] _result_T_212 = 8'h14 == de_bus_r_OP ? {{63'd0}, _result_T_79} : _result_T_210; // @[Mux.scala 81:58]
  wire [126:0] _result_T_214 = 8'h15 == de_bus_r_OP ? {{63'd0}, div_io_remainder} : _result_T_212; // @[Mux.scala 81:58]
  wire [126:0] _result_T_216 = 8'h16 == de_bus_r_OP ? {{63'd0}, div_io_remainder} : _result_T_214; // @[Mux.scala 81:58]
  wire [126:0] _result_T_218 = 8'h17 == de_bus_r_OP ? {{63'd0}, _result_T_84} : _result_T_216; // @[Mux.scala 81:58]
  wire [126:0] _result_T_220 = 8'h18 == de_bus_r_OP ? {{63'd0}, _result_T_84} : _result_T_218; // @[Mux.scala 81:58]
  wire [126:0] _result_T_222 = 8'h19 == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_220; // @[Mux.scala 81:58]
  wire [126:0] _result_T_224 = 8'h1a == de_bus_r_OP ? {{63'd0}, _result_T_99} : _result_T_222; // @[Mux.scala 81:58]
  wire [126:0] _result_T_226 = 8'h1b == de_bus_r_OP ? {{63'd0}, _result_T_101} : _result_T_224; // @[Mux.scala 81:58]
  wire [126:0] _result_T_228 = 8'h1c == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_226; // @[Mux.scala 81:58]
  wire [126:0] _result_T_230 = 8'h1d == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_228; // @[Mux.scala 81:58]
  wire [126:0] _result_T_232 = 8'h1e == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_230; // @[Mux.scala 81:58]
  wire [126:0] _result_T_234 = 8'h1f == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_232; // @[Mux.scala 81:58]
  wire [126:0] _result_T_236 = 8'h21 == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_234; // @[Mux.scala 81:58]
  wire [126:0] _result_T_238 = 8'h22 == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_236; // @[Mux.scala 81:58]
  wire [126:0] _result_T_240 = 8'h20 == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_238; // @[Mux.scala 81:58]
  wire [126:0] _result_T_242 = 8'h23 == de_bus_r_OP ? _result_T_117 : _result_T_240; // @[Mux.scala 81:58]
  wire [126:0] _result_T_244 = 8'h24 == de_bus_r_OP ? {{63'd0}, _result_T_125} : _result_T_242; // @[Mux.scala 81:58]
  wire [126:0] _result_T_246 = 8'h25 == de_bus_r_OP ? {{63'd0}, _result_T_127} : _result_T_244; // @[Mux.scala 81:58]
  wire [126:0] _result_T_248 = 8'h26 == de_bus_r_OP ? {{63'd0}, _result_T_135} : _result_T_246; // @[Mux.scala 81:58]
  wire [126:0] _result_T_250 = 8'h29 == de_bus_r_OP ? {{126'd0}, _result_T_138} : _result_T_248; // @[Mux.scala 81:58]
  wire [126:0] _result_T_252 = 8'h2a == de_bus_r_OP ? {{126'd0}, _result_T_140} : _result_T_250; // @[Mux.scala 81:58]
  wire [126:0] _result_T_254 = 8'h2b == de_bus_r_OP ? {{63'd0}, _result_T_142} : _result_T_252; // @[Mux.scala 81:58]
  wire [126:0] _result_T_256 = 8'h2c == de_bus_r_OP ? {{63'd0}, _result_T_143} : _result_T_254; // @[Mux.scala 81:58]
  wire [126:0] _result_T_258 = 8'h2d == de_bus_r_OP ? {{63'd0}, _result_T_144} : _result_T_256; // @[Mux.scala 81:58]
  wire [126:0] _result_T_260 = 8'h27 == de_bus_r_OP ? {{63'd0}, _result_T_148} : _result_T_258; // @[Mux.scala 81:58]
  wire [126:0] _result_T_262 = 8'h28 == de_bus_r_OP ? {{63'd0}, _result_T_158} : _result_T_260; // @[Mux.scala 81:58]
  wire [126:0] _result_T_264 = 8'h3c == de_bus_r_OP ? {{63'd0}, de_bus_r_csr_rdata} : _result_T_262; // @[Mux.scala 81:58]
  wire [126:0] _result_T_266 = 8'h3d == de_bus_r_OP ? {{63'd0}, de_bus_r_csr_rdata} : _result_T_264; // @[Mux.scala 81:58]
  wire [126:0] _result_T_268 = 8'h3e == de_bus_r_OP ? {{63'd0}, de_bus_r_csr_rdata} : _result_T_266; // @[Mux.scala 81:58]
  wire [126:0] _result_T_270 = 8'h2e == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_268; // @[Mux.scala 81:58]
  wire [126:0] _result_T_272 = 8'h31 == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_270; // @[Mux.scala 81:58]
  wire [126:0] _result_T_274 = 8'h30 == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_272; // @[Mux.scala 81:58]
  wire [126:0] _result_T_276 = 8'h2f == de_bus_r_OP ? {{63'd0}, _result_T_91} : _result_T_274; // @[Mux.scala 81:58]
  wire [126:0] _result_T_278 = 8'h38 == de_bus_r_OP ? {{63'd0}, de_bus_r_imm} : _result_T_276; // @[Mux.scala 81:58]
  wire [126:0] _result_T_280 = 8'h39 == de_bus_r_OP ? {{63'd0}, _result_T_168} : _result_T_278; // @[Mux.scala 81:58]
  wire [126:0] _result_T_282 = 8'h3a == de_bus_r_OP ? {{63'd0}, _result_T_101} : _result_T_280; // @[Mux.scala 81:58]
  wire [63:0] _csr_wdata_T = de_bus_r_csr_rdata | de_bus_r_rdata1; // @[EXU.scala 163:40]
  wire [63:0] _csr_wdata_T_1 = ~de_bus_r_rdata1; // @[EXU.scala 164:42]
  wire [63:0] _csr_wdata_T_2 = de_bus_r_csr_rdata & _csr_wdata_T_1; // @[EXU.scala 164:40]
  wire [63:0] _csr_wdata_T_4 = 8'h3c == de_bus_r_OP ? de_bus_r_rdata1 : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] _csr_wdata_T_6 = 8'h3d == de_bus_r_OP ? _csr_wdata_T : _csr_wdata_T_4; // @[Mux.scala 81:58]
  wire [63:0] _csr_wdata_T_8 = 8'h3e == de_bus_r_OP ? _csr_wdata_T_2 : _csr_wdata_T_6; // @[Mux.scala 81:58]
  wire  mul_end = mul_io_out_valid | mul_1_io_out_valid; // @[EXU.scala 202:34]
  wire  muling = is_mul_64 & ~mul_io_out_valid | is_mul_32 & ~mul_1_io_out_valid; // @[EXU.scala 203:50]
  wire  div_end = div_io_out_valid | div_1_io_out_valid; // @[EXU.scala 204:34]
  wire  _diving_T = ~div_io_out_valid; // @[EXU.scala 205:31]
  wire  _diving_T_2 = ~div_1_io_out_valid; // @[EXU.scala 205:67]
  wire  diving = is_div_64 & ~div_io_out_valid | is_div_32 & ~div_1_io_out_valid; // @[EXU.scala 205:50]
  wire  reming = is_rem_64 & _diving_T | is_rem_32 & _diving_T_2; // @[EXU.scala 206:50]
  wire  _es_ready_go_T_3 = muling | diving | reming ? 1'h0 : 1'h1; // @[EXU.scala 208:27]
  wire  es_ready_go = mul_end | div_end | _es_ready_go_T_3; // @[EXU.scala 207:27]
  mul mul ( // @[EXU.scala 51:23]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_mul_valid(mul_io_mul_valid),
    .io_multiplicand(mul_io_multiplicand),
    .io_multiplier(mul_io_multiplier),
    .io_out_valid(mul_io_out_valid),
    .io_result_lo(mul_io_result_lo)
  );
  mul_1 mul_1 ( // @[EXU.scala 52:23]
    .clock(mul_1_clock),
    .reset(mul_1_reset),
    .io_mul_valid(mul_1_io_mul_valid),
    .io_multiplicand(mul_1_io_multiplicand),
    .io_multiplier(mul_1_io_multiplier),
    .io_out_valid(mul_1_io_out_valid),
    .io_result_lo(mul_1_io_result_lo)
  );
  div div ( // @[EXU.scala 70:23]
    .clock(div_clock),
    .reset(div_reset),
    .io_dividend(div_io_dividend),
    .io_divisor(div_io_divisor),
    .io_div_valid(div_io_div_valid),
    .io_div_signed(div_io_div_signed),
    .io_out_valid(div_io_out_valid),
    .io_quotient(div_io_quotient),
    .io_remainder(div_io_remainder)
  );
  div_1 div_1 ( // @[EXU.scala 71:23]
    .clock(div_1_clock),
    .reset(div_1_reset),
    .io_dividend(div_1_io_dividend),
    .io_divisor(div_1_io_divisor),
    .io_div_valid(div_1_io_div_valid),
    .io_div_signed(div_1_io_div_signed),
    .io_out_valid(div_1_io_out_valid),
    .io_quotient(div_1_io_quotient),
    .io_remainder(div_1_io_remainder)
  );
  assign io_es_allowin = ~es_valid | es_ready_go & io_ms_allowin; // @[EXU.scala 210:34]
  assign io_es_to_ms_valid = es_valid & es_ready_go; // @[EXU.scala 211:33]
  assign io_em_bus_res_from_mem = de_bus_r_res_from_mem; // @[EXU.scala 169:26]
  assign io_em_bus_gr_we = de_bus_r_gr_we; // @[EXU.scala 170:26]
  assign io_em_bus_dest = de_bus_r_dest; // @[EXU.scala 171:26]
  assign io_em_bus_alu_result = _result_T_282[63:0]; // @[EXU.scala 173:26]
  assign io_em_bus_ex_pc = ex_pc[31:0]; // @[EXU.scala 172:26]
  assign io_em_bus_ld_type = de_bus_r_ld_type; // @[EXU.scala 174:26]
  assign io_em_bus_inst = de_bus_r_inst; // @[EXU.scala 175:26]
  assign io_em_bus_csr_wdata = 8'h3f == de_bus_r_OP ? de_bus_r_rdata1 : _csr_wdata_T_8; // @[Mux.scala 81:58]
  assign io_em_bus_csr_wen = de_bus_r_csr_wen; // @[EXU.scala 178:26]
  assign io_em_bus_csr_waddr1 = de_bus_r_csr_waddr1; // @[EXU.scala 182:25]
  assign io_em_bus_csr_waddr2 = de_bus_r_csr_waddr2; // @[EXU.scala 183:25]
  assign io_em_bus_eval = de_bus_r_eval; // @[EXU.scala 185:24]
  assign io_em_bus_is_ld = de_bus_r_is_ld; // @[EXU.scala 188:25]
  assign io_em_bus_MemWen = de_bus_r_MemWen; // @[EXU.scala 190:24]
  assign io_em_bus_Memwdata = de_bus_r_rdata2; // @[EXU.scala 191:24]
  assign io_em_bus_wmask = de_bus_r_wmask; // @[EXU.scala 192:23]
  assign io_es_dest_valid_gr_we = de_bus_r_gr_we; // @[EXU.scala 195:36]
  assign io_es_dest_valid_es_valid = es_valid; // @[EXU.scala 197:36]
  assign io_es_dest_valid_dest = de_bus_r_dest; // @[EXU.scala 196:36]
  assign io_es_dest_valid_es_forward_data = _result_T_282[63:0]; // @[EXU.scala 194:36]
  assign io_es_dest_valid_es_is_ld = de_bus_r_is_ld; // @[EXU.scala 198:36]
  assign io_es_dest_valid_es_ready_go = mul_end | div_end | _es_ready_go_T_3; // @[EXU.scala 207:27]
  assign io_es_dest_valid_es_to_ms_valid = io_es_to_ms_valid; // @[EXU.scala 200:36]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_mul_valid = is_mul_64 & es_valid; // @[EXU.scala 56:33]
  assign mul_io_multiplicand = de_bus_r_rdata1; // @[EXU.scala 60:23]
  assign mul_io_multiplier = de_bus_r_rdata2; // @[EXU.scala 61:21]
  assign mul_1_clock = clock;
  assign mul_1_reset = reset;
  assign mul_1_io_mul_valid = is_mul_32 & es_valid; // @[EXU.scala 63:33]
  assign mul_1_io_multiplicand = de_bus_r_rdata1[31:0]; // @[EXU.scala 67:30]
  assign mul_1_io_multiplier = de_bus_r_rdata2[31:0]; // @[EXU.scala 68:28]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_dividend = de_bus_r_rdata1; // @[EXU.scala 81:19]
  assign div_io_divisor = de_bus_r_rdata2; // @[EXU.scala 82:18]
  assign div_io_div_valid = (is_div_64 | is_rem_64) & es_valid; // @[EXU.scala 77:48]
  assign div_io_div_signed = _is_div_64_T | _is_rem_64_T; // @[EXU.scala 80:48]
  assign div_1_clock = clock;
  assign div_1_reset = reset;
  assign div_1_io_dividend = de_bus_r_rdata1[31:0]; // @[EXU.scala 88:26]
  assign div_1_io_divisor = de_bus_r_rdata2[31:0]; // @[EXU.scala 89:25]
  assign div_1_io_div_valid = (is_div_32 | is_rem_32) & es_valid; // @[EXU.scala 84:48]
  assign div_1_io_div_signed = _is_div_32_T | _is_rem_32_T; // @[EXU.scala 87:49]
  always @(posedge clock) begin
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_OP <= 8'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_OP <= io_de_bus_OP; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_res_from_mem <= 1'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_res_from_mem <= io_de_bus_res_from_mem; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_gr_we <= 1'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_gr_we <= io_de_bus_gr_we; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_MemWen <= 1'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_MemWen <= io_de_bus_MemWen; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_wmask <= 8'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_wmask <= io_de_bus_wmask; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_ds_pc <= 32'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_ds_pc <= io_de_bus_ds_pc; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_dest <= 5'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_dest <= io_de_bus_dest; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_imm <= 64'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_imm <= io_de_bus_imm; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_rdata1 <= 64'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_rdata1 <= io_de_bus_rdata1; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_rdata2 <= 64'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_rdata2 <= io_de_bus_rdata2; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_ld_type <= 3'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_ld_type <= io_de_bus_ld_type; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_inst <= 32'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_inst <= io_de_bus_inst; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_csr_rdata <= 64'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_csr_rdata <= io_de_bus_csr_rdata; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_csr_waddr1 <= 3'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_csr_waddr1 <= io_de_bus_csr_waddr1; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_csr_waddr2 <= 3'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_csr_waddr2 <= io_de_bus_csr_waddr2; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_csr_wen <= 1'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_csr_wen <= io_de_bus_csr_wen; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_eval <= 1'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_eval <= io_de_bus_eval; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 23:28]
      de_bus_r_is_ld <= 1'h0; // @[EXU.scala 23:28]
    end else if (io_ds_to_es_valid & io_es_allowin) begin // @[EXU.scala 31:44]
      de_bus_r_is_ld <= io_de_bus_is_ld; // @[EXU.scala 32:14]
    end
    if (reset) begin // @[EXU.scala 24:28]
      es_valid <= 1'h0; // @[EXU.scala 24:28]
    end else if (io_es_allowin) begin // @[EXU.scala 27:23]
      es_valid <= io_ds_to_es_valid; // @[EXU.scala 28:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  de_bus_r_OP = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  de_bus_r_res_from_mem = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  de_bus_r_gr_we = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  de_bus_r_MemWen = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  de_bus_r_wmask = _RAND_4[7:0];
  _RAND_5 = {1{`RANDOM}};
  de_bus_r_ds_pc = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  de_bus_r_dest = _RAND_6[4:0];
  _RAND_7 = {2{`RANDOM}};
  de_bus_r_imm = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  de_bus_r_rdata1 = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  de_bus_r_rdata2 = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  de_bus_r_ld_type = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  de_bus_r_inst = _RAND_11[31:0];
  _RAND_12 = {2{`RANDOM}};
  de_bus_r_csr_rdata = _RAND_12[63:0];
  _RAND_13 = {1{`RANDOM}};
  de_bus_r_csr_waddr1 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  de_bus_r_csr_waddr2 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  de_bus_r_csr_wen = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  de_bus_r_eval = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  de_bus_r_is_ld = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  es_valid = _RAND_18[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MEM(
  input         clock,
  input         reset,
  output        io_ms_allowin,
  input         io_es_to_ms_valid,
  output        io_ms_to_ws_valid,
  input         io_em_bus_res_from_mem,
  input         io_em_bus_gr_we,
  input  [4:0]  io_em_bus_dest,
  input  [63:0] io_em_bus_alu_result,
  input  [31:0] io_em_bus_ex_pc,
  input  [2:0]  io_em_bus_ld_type,
  input  [31:0] io_em_bus_inst,
  input  [63:0] io_em_bus_csr_wdata,
  input         io_em_bus_csr_wen,
  input  [2:0]  io_em_bus_csr_waddr1,
  input  [2:0]  io_em_bus_csr_waddr2,
  input         io_em_bus_eval,
  input         io_em_bus_is_ld,
  input         io_em_bus_MemWen,
  input  [63:0] io_em_bus_Memwdata,
  input  [7:0]  io_em_bus_wmask,
  output        io_mw_bus_gr_we,
  output [4:0]  io_mw_bus_dest,
  output [63:0] io_mw_bus_final_result,
  output [31:0] io_mw_bus_mem_pc,
  output [31:0] io_mw_bus_inst,
  output [63:0] io_mw_bus_csr_wdata,
  output        io_mw_bus_csr_wen,
  output [2:0]  io_mw_bus_csr_waddr1,
  output [2:0]  io_mw_bus_csr_waddr2,
  output        io_mw_bus_eval,
  output        io_ms_dest_valid_gr_we,
  output        io_ms_dest_valid_ms_valid,
  output [4:0]  io_ms_dest_valid_dest,
  output [63:0] io_ms_dest_valid_ms_forward_data,
  output        io_ms_dest_valid_ms_is_ld,
  output        io_ms_dest_valid_ms_to_ws_valid,
  output        io_ms_dest_valid_ms_ready_go,
  input  [63:0] io_data_sram_rdata,
  output [63:0] io_mem_result,
  output [2:0]  io_ld_type,
  input         io_data_sram_data_ok,
  output        io_data_sram_req,
  output        io_data_sram_we,
  output [31:0] io_data_sram_addr,
  output [63:0] io_data_sram_wdata,
  output [7:0]  io_data_sram_wmask,
  input         io_data_sram_addr_ok
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  reg  ms_valid; // @[MEM.scala 31:28]
  reg  em_bus_r_res_from_mem; // @[MEM.scala 33:28]
  reg  em_bus_r_gr_we; // @[MEM.scala 33:28]
  reg [4:0] em_bus_r_dest; // @[MEM.scala 33:28]
  reg [63:0] em_bus_r_alu_result; // @[MEM.scala 33:28]
  reg [31:0] em_bus_r_ex_pc; // @[MEM.scala 33:28]
  reg [2:0] em_bus_r_ld_type; // @[MEM.scala 33:28]
  reg [31:0] em_bus_r_inst; // @[MEM.scala 33:28]
  reg [63:0] em_bus_r_csr_wdata; // @[MEM.scala 33:28]
  reg  em_bus_r_csr_wen; // @[MEM.scala 33:28]
  reg [2:0] em_bus_r_csr_waddr1; // @[MEM.scala 33:28]
  reg [2:0] em_bus_r_csr_waddr2; // @[MEM.scala 33:28]
  reg  em_bus_r_eval; // @[MEM.scala 33:28]
  reg  em_bus_r_is_ld; // @[MEM.scala 33:28]
  reg  em_bus_r_MemWen; // @[MEM.scala 33:28]
  reg [63:0] em_bus_r_Memwdata; // @[MEM.scala 33:28]
  reg [7:0] em_bus_r_wmask; // @[MEM.scala 33:28]
  reg  mid_handshake_data; // @[MEM.scala 35:37]
  wire  _ms_ready_go_T = em_bus_r_res_from_mem | em_bus_r_MemWen; // @[MEM.scala 37:50]
  wire  ms_ready_go = em_bus_r_res_from_mem | em_bus_r_MemWen ? io_data_sram_data_ok : 1'h1; // @[MEM.scala 37:27]
  wire  _GEN_62 = io_ms_allowin ? 1'h0 : mid_handshake_data; // @[MEM.scala 72:28 73:24 35:37]
  wire  _GEN_63 = io_data_sram_addr_ok & io_data_sram_req & ~io_ms_allowin | _GEN_62; // @[MEM.scala 70:73 71:24]
  wire [55:0] _io_mem_result_T_3 = io_data_sram_rdata[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_mem_result_T_4 = {_io_mem_result_T_3,io_data_sram_rdata[7:0]}; // @[Cat.scala 31:58]
  wire [47:0] _io_mem_result_T_8 = io_data_sram_rdata[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_mem_result_T_9 = {_io_mem_result_T_8,io_data_sram_rdata[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] _io_mem_result_T_13 = io_data_sram_rdata[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 74:12]
  wire [63:0] _io_mem_result_T_14 = {_io_mem_result_T_13,io_data_sram_rdata[31:0]}; // @[Cat.scala 31:58]
  wire [63:0] _io_mem_result_T_20 = 3'h0 == io_ld_type ? _io_mem_result_T_4 : io_data_sram_rdata; // @[Mux.scala 81:58]
  wire [63:0] _io_mem_result_T_22 = 3'h1 == io_ld_type ? _io_mem_result_T_9 : _io_mem_result_T_20; // @[Mux.scala 81:58]
  wire [63:0] _io_mem_result_T_24 = 3'h2 == io_ld_type ? _io_mem_result_T_14 : _io_mem_result_T_22; // @[Mux.scala 81:58]
  wire [63:0] _io_mem_result_T_26 = 3'h3 == io_ld_type ? io_data_sram_rdata : _io_mem_result_T_24; // @[Mux.scala 81:58]
  wire [63:0] _io_mem_result_T_28 = 3'h4 == io_ld_type ? {{56'd0}, io_data_sram_rdata[7:0]} : _io_mem_result_T_26; // @[Mux.scala 81:58]
  wire [63:0] _io_mem_result_T_30 = 3'h5 == io_ld_type ? {{48'd0}, io_data_sram_rdata[15:0]} : _io_mem_result_T_28; // @[Mux.scala 81:58]
  assign io_ms_allowin = ~ms_valid | ms_ready_go; // @[MEM.scala 38:34]
  assign io_ms_to_ws_valid = ms_valid & ms_ready_go; // @[MEM.scala 39:33]
  assign io_mw_bus_gr_we = em_bus_r_gr_we; // @[MEM.scala 103:26]
  assign io_mw_bus_dest = em_bus_r_dest; // @[MEM.scala 104:26]
  assign io_mw_bus_final_result = em_bus_r_res_from_mem ? io_mem_result : em_bus_r_alu_result; // @[MEM.scala 93:42]
  assign io_mw_bus_mem_pc = em_bus_r_ex_pc; // @[MEM.scala 106:26]
  assign io_mw_bus_inst = em_bus_r_inst; // @[MEM.scala 107:26]
  assign io_mw_bus_csr_wdata = em_bus_r_csr_wdata; // @[MEM.scala 109:26]
  assign io_mw_bus_csr_wen = em_bus_r_csr_wen; // @[MEM.scala 110:26]
  assign io_mw_bus_csr_waddr1 = em_bus_r_csr_waddr1; // @[MEM.scala 111:26]
  assign io_mw_bus_csr_waddr2 = em_bus_r_csr_waddr2; // @[MEM.scala 112:26]
  assign io_mw_bus_eval = em_bus_r_eval; // @[MEM.scala 115:26]
  assign io_ms_dest_valid_gr_we = em_bus_r_gr_we; // @[MEM.scala 96:29]
  assign io_ms_dest_valid_ms_valid = ms_valid; // @[MEM.scala 98:29]
  assign io_ms_dest_valid_dest = em_bus_r_dest; // @[MEM.scala 97:29]
  assign io_ms_dest_valid_ms_forward_data = em_bus_r_res_from_mem ? io_mem_result : em_bus_r_alu_result; // @[MEM.scala 93:42]
  assign io_ms_dest_valid_ms_is_ld = em_bus_r_is_ld; // @[MEM.scala 99:29]
  assign io_ms_dest_valid_ms_to_ws_valid = io_ms_to_ws_valid; // @[MEM.scala 100:35]
  assign io_ms_dest_valid_ms_ready_go = em_bus_r_res_from_mem | em_bus_r_MemWen ? io_data_sram_data_ok : 1'h1; // @[MEM.scala 37:27]
  assign io_mem_result = 3'h6 == io_ld_type ? {{32'd0}, io_data_sram_rdata[31:0]} : _io_mem_result_T_30; // @[Mux.scala 81:58]
  assign io_ld_type = em_bus_r_ld_type; // @[MEM.scala 120:26]
  assign io_data_sram_req = _ms_ready_go_T & ~mid_handshake_data & ms_valid; // @[MEM.scala 127:91]
  assign io_data_sram_we = em_bus_r_MemWen; // @[MEM.scala 123:22]
  assign io_data_sram_addr = em_bus_r_alu_result[31:0]; // @[MEM.scala 124:22]
  assign io_data_sram_wdata = em_bus_r_Memwdata; // @[MEM.scala 125:22]
  assign io_data_sram_wmask = em_bus_r_wmask; // @[MEM.scala 126:22]
  always @(posedge clock) begin
    if (reset) begin // @[MEM.scala 31:28]
      ms_valid <= 1'h0; // @[MEM.scala 31:28]
    end else if (io_ms_allowin) begin // @[MEM.scala 41:23]
      ms_valid <= io_es_to_ms_valid; // @[MEM.scala 42:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_res_from_mem <= 1'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_res_from_mem <= io_em_bus_res_from_mem; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_gr_we <= 1'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_gr_we <= io_em_bus_gr_we; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_dest <= 5'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_dest <= io_em_bus_dest; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_alu_result <= 64'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_alu_result <= io_em_bus_alu_result; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_ex_pc <= 32'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_ex_pc <= io_em_bus_ex_pc; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_ld_type <= 3'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_ld_type <= io_em_bus_ld_type; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_inst <= 32'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_inst <= io_em_bus_inst; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_csr_wdata <= 64'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_csr_wdata <= io_em_bus_csr_wdata; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_csr_wen <= 1'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_csr_wen <= io_em_bus_csr_wen; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_csr_waddr1 <= 3'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_csr_waddr1 <= io_em_bus_csr_waddr1; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_csr_waddr2 <= 3'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_csr_waddr2 <= io_em_bus_csr_waddr2; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_eval <= 1'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_eval <= io_em_bus_eval; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_is_ld <= 1'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_is_ld <= io_em_bus_is_ld; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_MemWen <= 1'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_MemWen <= io_em_bus_MemWen; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_Memwdata <= 64'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_Memwdata <= io_em_bus_Memwdata; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 33:28]
      em_bus_r_wmask <= 8'h0; // @[MEM.scala 33:28]
    end else if (io_es_to_ms_valid & io_ms_allowin) begin // @[MEM.scala 45:44]
      em_bus_r_wmask <= io_em_bus_wmask; // @[MEM.scala 46:14]
    end
    if (reset) begin // @[MEM.scala 35:37]
      mid_handshake_data <= 1'h0; // @[MEM.scala 35:37]
    end else if (io_data_sram_data_ok) begin // @[MEM.scala 68:29]
      mid_handshake_data <= 1'h0; // @[MEM.scala 69:24]
    end else begin
      mid_handshake_data <= _GEN_63;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ms_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  em_bus_r_res_from_mem = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  em_bus_r_gr_we = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  em_bus_r_dest = _RAND_3[4:0];
  _RAND_4 = {2{`RANDOM}};
  em_bus_r_alu_result = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  em_bus_r_ex_pc = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  em_bus_r_ld_type = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  em_bus_r_inst = _RAND_7[31:0];
  _RAND_8 = {2{`RANDOM}};
  em_bus_r_csr_wdata = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  em_bus_r_csr_wen = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  em_bus_r_csr_waddr1 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  em_bus_r_csr_waddr2 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  em_bus_r_eval = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  em_bus_r_is_ld = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  em_bus_r_MemWen = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  em_bus_r_Memwdata = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  em_bus_r_wmask = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  mid_handshake_data = _RAND_17[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module WBU(
  input         clock,
  input         reset,
  output        io_ws_allowin,
  input         io_ms_to_ws_valid,
  input         io_mw_bus_gr_we,
  input  [4:0]  io_mw_bus_dest,
  input  [63:0] io_mw_bus_final_result,
  input  [31:0] io_mw_bus_mem_pc,
  input  [31:0] io_mw_bus_inst,
  input  [63:0] io_mw_bus_csr_wdata,
  input         io_mw_bus_csr_wen,
  input  [2:0]  io_mw_bus_csr_waddr1,
  input  [2:0]  io_mw_bus_csr_waddr2,
  input         io_mw_bus_eval,
  output        io_rf_bus_rf_we,
  output [4:0]  io_rf_bus_rf_waddr,
  output [63:0] io_rf_bus_rf_wdata,
  output [31:0] io_rf_bus_wb_pc,
  output [31:0] io_rf_bus_wb_inst,
  output [63:0] io_rf_bus_csr_wdata,
  output        io_rf_bus_csr_wen,
  output [2:0]  io_rf_bus_csr_waddr1,
  output [2:0]  io_rf_bus_csr_waddr2,
  output        io_rf_bus_eval,
  output        io_in_WB,
  output        io_ws_dest_valid_gr_we,
  output        io_ws_dest_valid_ws_valid,
  output [4:0]  io_ws_dest_valid_dest,
  output [63:0] io_ws_dest_valid_ws_forward_data,
  output [63:0] io_wb_pc,
  output [63:0] io_wb_inst
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg  ws_valid; // @[WBU.scala 21:28]
  reg  mw_bus_r_gr_we; // @[WBU.scala 22:28]
  reg [4:0] mw_bus_r_dest; // @[WBU.scala 22:28]
  reg [63:0] mw_bus_r_final_result; // @[WBU.scala 22:28]
  reg [31:0] mw_bus_r_mem_pc; // @[WBU.scala 22:28]
  reg [31:0] mw_bus_r_inst; // @[WBU.scala 22:28]
  reg [63:0] mw_bus_r_csr_wdata; // @[WBU.scala 22:28]
  reg  mw_bus_r_csr_wen; // @[WBU.scala 22:28]
  reg [2:0] mw_bus_r_csr_waddr1; // @[WBU.scala 22:28]
  reg [2:0] mw_bus_r_csr_waddr2; // @[WBU.scala 22:28]
  reg  mw_bus_r_eval; // @[WBU.scala 22:28]
  assign io_ws_allowin = 1'h1; // @[WBU.scala 25:30]
  assign io_rf_bus_rf_we = mw_bus_r_gr_we & ws_valid; // @[WBU.scala 45:30]
  assign io_rf_bus_rf_waddr = mw_bus_r_dest; // @[WBU.scala 50:22]
  assign io_rf_bus_rf_wdata = mw_bus_r_final_result; // @[WBU.scala 51:22]
  assign io_rf_bus_wb_pc = mw_bus_r_mem_pc; // @[WBU.scala 52:21]
  assign io_rf_bus_wb_inst = mw_bus_r_inst; // @[WBU.scala 53:21]
  assign io_rf_bus_csr_wdata = mw_bus_r_csr_wdata; // @[WBU.scala 57:23]
  assign io_rf_bus_csr_wen = mw_bus_r_csr_wen; // @[WBU.scala 58:21]
  assign io_rf_bus_csr_waddr1 = mw_bus_r_csr_waddr1; // @[WBU.scala 60:24]
  assign io_rf_bus_csr_waddr2 = mw_bus_r_csr_waddr2; // @[WBU.scala 61:24]
  assign io_rf_bus_eval = mw_bus_r_eval; // @[WBU.scala 54:21]
  assign io_in_WB = ws_valid; // @[WBU.scala 26:17]
  assign io_ws_dest_valid_gr_we = mw_bus_r_gr_we; // @[WBU.scala 72:36]
  assign io_ws_dest_valid_ws_valid = ws_valid; // @[WBU.scala 71:36]
  assign io_ws_dest_valid_dest = mw_bus_r_dest; // @[WBU.scala 73:36]
  assign io_ws_dest_valid_ws_forward_data = mw_bus_r_final_result; // @[WBU.scala 74:36]
  assign io_wb_pc = {{32'd0}, mw_bus_r_mem_pc}; // @[WBU.scala 55:22]
  assign io_wb_inst = {{32'd0}, mw_bus_r_inst}; // @[WBU.scala 56:22]
  always @(posedge clock) begin
    if (reset) begin // @[WBU.scala 21:28]
      ws_valid <= 1'h0; // @[WBU.scala 21:28]
    end else if (io_ws_allowin) begin // @[WBU.scala 34:23]
      ws_valid <= io_ms_to_ws_valid; // @[WBU.scala 35:14]
    end
    if (reset) begin // @[WBU.scala 22:28]
      mw_bus_r_gr_we <= 1'h0; // @[WBU.scala 22:28]
    end else if (io_ms_to_ws_valid & io_ws_allowin) begin // @[WBU.scala 38:44]
      mw_bus_r_gr_we <= io_mw_bus_gr_we; // @[WBU.scala 39:14]
    end
    if (reset) begin // @[WBU.scala 22:28]
      mw_bus_r_dest <= 5'h0; // @[WBU.scala 22:28]
    end else if (io_ms_to_ws_valid & io_ws_allowin) begin // @[WBU.scala 38:44]
      mw_bus_r_dest <= io_mw_bus_dest; // @[WBU.scala 39:14]
    end
    if (reset) begin // @[WBU.scala 22:28]
      mw_bus_r_final_result <= 64'h0; // @[WBU.scala 22:28]
    end else if (io_ms_to_ws_valid & io_ws_allowin) begin // @[WBU.scala 38:44]
      mw_bus_r_final_result <= io_mw_bus_final_result; // @[WBU.scala 39:14]
    end
    if (reset) begin // @[WBU.scala 22:28]
      mw_bus_r_mem_pc <= 32'h0; // @[WBU.scala 22:28]
    end else if (io_ms_to_ws_valid & io_ws_allowin) begin // @[WBU.scala 38:44]
      mw_bus_r_mem_pc <= io_mw_bus_mem_pc; // @[WBU.scala 39:14]
    end
    if (reset) begin // @[WBU.scala 22:28]
      mw_bus_r_inst <= 32'h0; // @[WBU.scala 22:28]
    end else if (io_ms_to_ws_valid & io_ws_allowin) begin // @[WBU.scala 38:44]
      mw_bus_r_inst <= io_mw_bus_inst; // @[WBU.scala 39:14]
    end
    if (reset) begin // @[WBU.scala 22:28]
      mw_bus_r_csr_wdata <= 64'h0; // @[WBU.scala 22:28]
    end else if (io_ms_to_ws_valid & io_ws_allowin) begin // @[WBU.scala 38:44]
      mw_bus_r_csr_wdata <= io_mw_bus_csr_wdata; // @[WBU.scala 39:14]
    end
    if (reset) begin // @[WBU.scala 22:28]
      mw_bus_r_csr_wen <= 1'h0; // @[WBU.scala 22:28]
    end else if (io_ms_to_ws_valid & io_ws_allowin) begin // @[WBU.scala 38:44]
      mw_bus_r_csr_wen <= io_mw_bus_csr_wen; // @[WBU.scala 39:14]
    end
    if (reset) begin // @[WBU.scala 22:28]
      mw_bus_r_csr_waddr1 <= 3'h0; // @[WBU.scala 22:28]
    end else if (io_ms_to_ws_valid & io_ws_allowin) begin // @[WBU.scala 38:44]
      mw_bus_r_csr_waddr1 <= io_mw_bus_csr_waddr1; // @[WBU.scala 39:14]
    end
    if (reset) begin // @[WBU.scala 22:28]
      mw_bus_r_csr_waddr2 <= 3'h0; // @[WBU.scala 22:28]
    end else if (io_ms_to_ws_valid & io_ws_allowin) begin // @[WBU.scala 38:44]
      mw_bus_r_csr_waddr2 <= io_mw_bus_csr_waddr2; // @[WBU.scala 39:14]
    end
    if (reset) begin // @[WBU.scala 22:28]
      mw_bus_r_eval <= 1'h0; // @[WBU.scala 22:28]
    end else if (io_ms_to_ws_valid & io_ws_allowin) begin // @[WBU.scala 38:44]
      mw_bus_r_eval <= io_mw_bus_eval; // @[WBU.scala 39:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ws_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  mw_bus_r_gr_we = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mw_bus_r_dest = _RAND_2[4:0];
  _RAND_3 = {2{`RANDOM}};
  mw_bus_r_final_result = _RAND_3[63:0];
  _RAND_4 = {1{`RANDOM}};
  mw_bus_r_mem_pc = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  mw_bus_r_inst = _RAND_5[31:0];
  _RAND_6 = {2{`RANDOM}};
  mw_bus_r_csr_wdata = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  mw_bus_r_csr_wen = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  mw_bus_r_csr_waddr1 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  mw_bus_r_csr_waddr2 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  mw_bus_r_eval = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AXI(
  input          clock,
  input          reset,
  output [3:0]   io_arid,
  output [63:0]  io_araddr,
  output         io_arvalid,
  input          io_arready,
  input  [63:0]  io_rdata,
  input  [127:0] io_icache_rdata,
  input          io_rvalid,
  output         io_rready,
  output [63:0]  io_awaddr,
  output         io_awvalid,
  input          io_awready,
  output [63:0]  io_wdata,
  output [7:0]   io_wstrb,
  output         io_wvalid,
  input          io_wready,
  input          io_bvalid,
  output         io_bready,
  input          io_inst_sram_req,
  input  [63:0]  io_inst_sram_addr,
  output [127:0] io_inst_sram_rdata,
  output         io_inst_sram_addr_ok,
  output         io_inst_sram_data_ok,
  input          io_data_sram_req,
  input          io_data_sram_wr,
  input  [7:0]   io_data_sram_wstrb,
  input  [63:0]  io_data_sram_addr,
  input  [63:0]  io_data_sram_wdata,
  output [63:0]  io_data_sram_rdata,
  output         io_data_sram_addr_ok,
  output         io_data_sram_data_ok
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] rstate; // @[AXI.scala 72:55]
  wire  read_ainit = rstate == 2'h0; // @[AXI.scala 74:29]
  wire  read_araddr = rstate == 2'h1; // @[AXI.scala 75:29]
  wire  read_rdata = rstate == 2'h2; // @[AXI.scala 76:29]
  reg  reading_inst_sram; // @[AXI.scala 78:34]
  reg  reading_data_sram; // @[AXI.scala 79:34]
  reg [1:0] wstate; // @[AXI.scala 85:76]
  wire  write_init = wstate == 2'h0; // @[AXI.scala 87:28]
  wire  write_addr = wstate == 2'h1; // @[AXI.scala 88:28]
  wire  write_data = wstate == 2'h2; // @[AXI.scala 89:28]
  reg [1:0] writing_data_sram; // @[AXI.scala 92:34]
  wire  _T_2 = io_data_sram_req & ~io_data_sram_wr; // @[AXI.scala 96:31]
  wire [1:0] _GEN_2 = io_rvalid ? 2'h0 : 2'h2; // @[AXI.scala 110:23 111:16 113:16]
  wire  _T_16 = read_rdata & io_rvalid & io_rready; // @[AXI.scala 121:38]
  wire  _GEN_6 = read_rdata & io_rvalid & io_rready ? 1'h0 : reading_inst_sram; // @[AXI.scala 121:52 122:23 124:23]
  wire  _GEN_7 = ~io_data_sram_req & io_inst_sram_req & write_init & read_ainit | _GEN_6; // @[AXI.scala 119:95 120:23]
  wire  _GEN_8 = _T_16 ? 1'h0 : reading_data_sram; // @[AXI.scala 130:52 131:23 79:34]
  wire  _GEN_9 = _T_2 & write_init & read_ainit | _GEN_8; // @[AXI.scala 128:74 129:23]
  wire  _io_arid_T = read_araddr & reading_data_sram; // @[AXI.scala 135:33]
  wire  _io_arid_T_1 = read_araddr & reading_inst_sram; // @[AXI.scala 135:76]
  wire [1:0] _io_arid_T_2 = read_araddr & reading_inst_sram ? 2'h0 : 2'h2; // @[AXI.scala 135:63]
  wire [1:0] _io_arid_T_3 = read_araddr & reading_data_sram ? 2'h1 : _io_arid_T_2; // @[AXI.scala 135:20]
  wire [63:0] _io_araddr_T_2 = _io_arid_T_1 ? io_inst_sram_addr : 64'h0; // @[AXI.scala 140:8]
  wire [1:0] _GEN_12 = io_wready ? 2'h3 : 2'h2; // @[AXI.scala 161:23 162:16 164:16]
  wire [1:0] _GEN_13 = io_bvalid ? 2'h0 : wstate; // @[AXI.scala 168:23 169:16 85:76]
  wire [1:0] _GEN_14 = 2'h3 == wstate ? _GEN_13 : wstate; // @[AXI.scala 145:18 85:76]
  wire [1:0] _writing_data_sram_T_1 = writing_data_sram + 2'h1; // @[AXI.scala 178:44]
  assign io_arid = {{2'd0}, _io_arid_T_3}; // @[AXI.scala 135:14]
  assign io_araddr = _io_arid_T ? io_data_sram_addr : _io_araddr_T_2; // @[AXI.scala 137:19]
  assign io_arvalid = rstate == 2'h1; // @[AXI.scala 75:29]
  assign io_rready = rstate == 2'h2; // @[AXI.scala 76:29]
  assign io_awaddr = write_addr ? io_data_sram_addr : 64'h0; // @[AXI.scala 184:20]
  assign io_awvalid = wstate == 2'h1; // @[AXI.scala 88:28]
  assign io_wdata = write_data ? io_data_sram_wdata : 64'h0; // @[AXI.scala 187:19]
  assign io_wstrb = write_data ? io_data_sram_wstrb : 8'h0; // @[AXI.scala 188:19]
  assign io_wvalid = wstate == 2'h2; // @[AXI.scala 89:28]
  assign io_bready = wstate == 2'h3; // @[AXI.scala 90:28]
  assign io_inst_sram_rdata = io_icache_rdata; // @[AXI.scala 197:24]
  assign io_inst_sram_addr_ok = reading_inst_sram & io_arready; // @[AXI.scala 192:45]
  assign io_inst_sram_data_ok = reading_inst_sram & io_rvalid; // @[AXI.scala 194:45]
  assign io_data_sram_rdata = io_rdata; // @[AXI.scala 196:24]
  assign io_data_sram_addr_ok = reading_data_sram & io_arready | writing_data_sram == 2'h2; // @[AXI.scala 193:59]
  assign io_data_sram_data_ok = reading_data_sram & io_rvalid | io_bready; // @[AXI.scala 195:58]
  always @(posedge clock) begin
    if (reset) begin // @[AXI.scala 72:55]
      rstate <= 2'h0; // @[AXI.scala 72:55]
    end else if (2'h0 == rstate) begin // @[AXI.scala 94:18]
      if ((io_data_sram_req & ~io_data_sram_wr | io_inst_sram_req) & write_init) begin // @[AXI.scala 96:110]
        rstate <= 2'h1; // @[AXI.scala 97:16]
      end else begin
        rstate <= 2'h0; // @[AXI.scala 99:16]
      end
    end else if (2'h1 == rstate) begin // @[AXI.scala 94:18]
      if (io_arready) begin // @[AXI.scala 103:24]
        rstate <= 2'h2; // @[AXI.scala 104:16]
      end else begin
        rstate <= 2'h1; // @[AXI.scala 106:16]
      end
    end else if (2'h2 == rstate) begin // @[AXI.scala 94:18]
      rstate <= _GEN_2;
    end
    if (reset) begin // @[AXI.scala 78:34]
      reading_inst_sram <= 1'h0; // @[AXI.scala 78:34]
    end else begin
      reading_inst_sram <= _GEN_7;
    end
    if (reset) begin // @[AXI.scala 79:34]
      reading_data_sram <= 1'h0; // @[AXI.scala 79:34]
    end else begin
      reading_data_sram <= _GEN_9;
    end
    if (reset) begin // @[AXI.scala 85:76]
      wstate <= 2'h0; // @[AXI.scala 85:76]
    end else if (2'h0 == wstate) begin // @[AXI.scala 145:18]
      if (io_data_sram_req & io_data_sram_wr) begin // @[AXI.scala 147:51]
        wstate <= 2'h1; // @[AXI.scala 148:16]
      end else begin
        wstate <= 2'h0; // @[AXI.scala 150:16]
      end
    end else if (2'h1 == wstate) begin // @[AXI.scala 145:18]
      if (io_awready) begin // @[AXI.scala 154:24]
        wstate <= 2'h2; // @[AXI.scala 155:16]
      end else begin
        wstate <= 2'h1; // @[AXI.scala 157:16]
      end
    end else if (2'h2 == wstate) begin // @[AXI.scala 145:18]
      wstate <= _GEN_12;
    end else begin
      wstate <= _GEN_14;
    end
    if (reset) begin // @[AXI.scala 92:34]
      writing_data_sram <= 2'h0; // @[AXI.scala 92:34]
    end else if (io_awready | io_wready) begin // @[AXI.scala 177:39]
      writing_data_sram <= _writing_data_sram_T_1; // @[AXI.scala 178:23]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rstate = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  reading_inst_sram = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  reading_data_sram = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  wstate = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  writing_data_sram = _RAND_4[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module icache(
  input          clock,
  input          reset,
  input          io_valid,
  input  [63:0]  io_addr,
  output [63:0]  io_rdata,
  output         io_addr_ok,
  output         io_data_ok,
  output         io_rd_req,
  output [31:0]  io_rd_addr,
  input          io_rd_rdy,
  input  [127:0] io_rd_data,
  input          io_inst_sram_data_ok
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [191:0] _RAND_3;
  reg [191:0] _RAND_4;
  reg [191:0] _RAND_5;
  reg [191:0] _RAND_6;
  reg [191:0] _RAND_7;
  reg [191:0] _RAND_8;
  reg [191:0] _RAND_9;
  reg [191:0] _RAND_10;
  reg [191:0] _RAND_11;
  reg [191:0] _RAND_12;
  reg [191:0] _RAND_13;
  reg [191:0] _RAND_14;
  reg [191:0] _RAND_15;
  reg [191:0] _RAND_16;
  reg [191:0] _RAND_17;
  reg [191:0] _RAND_18;
  reg [191:0] _RAND_19;
  reg [191:0] _RAND_20;
  reg [191:0] _RAND_21;
  reg [191:0] _RAND_22;
  reg [191:0] _RAND_23;
  reg [191:0] _RAND_24;
  reg [191:0] _RAND_25;
  reg [191:0] _RAND_26;
  reg [191:0] _RAND_27;
  reg [191:0] _RAND_28;
  reg [191:0] _RAND_29;
  reg [191:0] _RAND_30;
  reg [191:0] _RAND_31;
  reg [191:0] _RAND_32;
  reg [191:0] _RAND_33;
  reg [191:0] _RAND_34;
  reg [191:0] _RAND_35;
  reg [191:0] _RAND_36;
  reg [191:0] _RAND_37;
  reg [191:0] _RAND_38;
  reg [191:0] _RAND_39;
  reg [191:0] _RAND_40;
  reg [191:0] _RAND_41;
  reg [191:0] _RAND_42;
  reg [191:0] _RAND_43;
  reg [191:0] _RAND_44;
  reg [191:0] _RAND_45;
  reg [191:0] _RAND_46;
  reg [191:0] _RAND_47;
  reg [191:0] _RAND_48;
  reg [191:0] _RAND_49;
  reg [191:0] _RAND_50;
  reg [191:0] _RAND_51;
  reg [191:0] _RAND_52;
  reg [191:0] _RAND_53;
  reg [191:0] _RAND_54;
  reg [191:0] _RAND_55;
  reg [191:0] _RAND_56;
  reg [191:0] _RAND_57;
  reg [191:0] _RAND_58;
  reg [191:0] _RAND_59;
  reg [191:0] _RAND_60;
  reg [191:0] _RAND_61;
  reg [191:0] _RAND_62;
  reg [191:0] _RAND_63;
  reg [191:0] _RAND_64;
  reg [191:0] _RAND_65;
  reg [191:0] _RAND_66;
  reg [191:0] _RAND_67;
  reg [191:0] _RAND_68;
  reg [191:0] _RAND_69;
  reg [191:0] _RAND_70;
  reg [191:0] _RAND_71;
  reg [191:0] _RAND_72;
  reg [191:0] _RAND_73;
  reg [191:0] _RAND_74;
  reg [191:0] _RAND_75;
  reg [191:0] _RAND_76;
  reg [191:0] _RAND_77;
  reg [191:0] _RAND_78;
  reg [191:0] _RAND_79;
  reg [191:0] _RAND_80;
  reg [191:0] _RAND_81;
  reg [191:0] _RAND_82;
  reg [191:0] _RAND_83;
  reg [191:0] _RAND_84;
  reg [191:0] _RAND_85;
  reg [191:0] _RAND_86;
  reg [191:0] _RAND_87;
  reg [191:0] _RAND_88;
  reg [191:0] _RAND_89;
  reg [191:0] _RAND_90;
  reg [191:0] _RAND_91;
  reg [191:0] _RAND_92;
  reg [191:0] _RAND_93;
  reg [191:0] _RAND_94;
  reg [191:0] _RAND_95;
  reg [191:0] _RAND_96;
  reg [191:0] _RAND_97;
  reg [191:0] _RAND_98;
  reg [191:0] _RAND_99;
  reg [191:0] _RAND_100;
  reg [191:0] _RAND_101;
  reg [191:0] _RAND_102;
  reg [191:0] _RAND_103;
  reg [191:0] _RAND_104;
  reg [191:0] _RAND_105;
  reg [191:0] _RAND_106;
  reg [191:0] _RAND_107;
  reg [191:0] _RAND_108;
  reg [191:0] _RAND_109;
  reg [191:0] _RAND_110;
  reg [191:0] _RAND_111;
  reg [191:0] _RAND_112;
  reg [191:0] _RAND_113;
  reg [191:0] _RAND_114;
  reg [191:0] _RAND_115;
  reg [191:0] _RAND_116;
  reg [191:0] _RAND_117;
  reg [191:0] _RAND_118;
  reg [191:0] _RAND_119;
  reg [191:0] _RAND_120;
  reg [191:0] _RAND_121;
  reg [191:0] _RAND_122;
  reg [191:0] _RAND_123;
  reg [191:0] _RAND_124;
  reg [191:0] _RAND_125;
  reg [191:0] _RAND_126;
  reg [191:0] _RAND_127;
  reg [191:0] _RAND_128;
  reg [191:0] _RAND_129;
  reg [191:0] _RAND_130;
  reg [191:0] _RAND_131;
  reg [191:0] _RAND_132;
  reg [191:0] _RAND_133;
  reg [191:0] _RAND_134;
  reg [191:0] _RAND_135;
  reg [191:0] _RAND_136;
  reg [191:0] _RAND_137;
  reg [191:0] _RAND_138;
  reg [191:0] _RAND_139;
  reg [191:0] _RAND_140;
  reg [191:0] _RAND_141;
  reg [191:0] _RAND_142;
  reg [191:0] _RAND_143;
  reg [191:0] _RAND_144;
  reg [191:0] _RAND_145;
  reg [191:0] _RAND_146;
  reg [191:0] _RAND_147;
  reg [191:0] _RAND_148;
  reg [191:0] _RAND_149;
  reg [191:0] _RAND_150;
  reg [191:0] _RAND_151;
  reg [191:0] _RAND_152;
  reg [191:0] _RAND_153;
  reg [191:0] _RAND_154;
  reg [191:0] _RAND_155;
  reg [191:0] _RAND_156;
  reg [191:0] _RAND_157;
  reg [191:0] _RAND_158;
  reg [191:0] _RAND_159;
  reg [191:0] _RAND_160;
  reg [191:0] _RAND_161;
  reg [191:0] _RAND_162;
  reg [191:0] _RAND_163;
  reg [191:0] _RAND_164;
  reg [191:0] _RAND_165;
  reg [191:0] _RAND_166;
  reg [191:0] _RAND_167;
  reg [191:0] _RAND_168;
  reg [191:0] _RAND_169;
  reg [191:0] _RAND_170;
  reg [191:0] _RAND_171;
  reg [191:0] _RAND_172;
  reg [191:0] _RAND_173;
  reg [191:0] _RAND_174;
  reg [191:0] _RAND_175;
  reg [191:0] _RAND_176;
  reg [191:0] _RAND_177;
  reg [191:0] _RAND_178;
  reg [191:0] _RAND_179;
  reg [191:0] _RAND_180;
  reg [191:0] _RAND_181;
  reg [191:0] _RAND_182;
  reg [191:0] _RAND_183;
  reg [191:0] _RAND_184;
  reg [191:0] _RAND_185;
  reg [191:0] _RAND_186;
  reg [191:0] _RAND_187;
  reg [191:0] _RAND_188;
  reg [191:0] _RAND_189;
  reg [191:0] _RAND_190;
  reg [191:0] _RAND_191;
  reg [191:0] _RAND_192;
  reg [191:0] _RAND_193;
  reg [191:0] _RAND_194;
  reg [191:0] _RAND_195;
  reg [191:0] _RAND_196;
  reg [191:0] _RAND_197;
  reg [191:0] _RAND_198;
  reg [191:0] _RAND_199;
  reg [191:0] _RAND_200;
  reg [191:0] _RAND_201;
  reg [191:0] _RAND_202;
  reg [191:0] _RAND_203;
  reg [191:0] _RAND_204;
  reg [191:0] _RAND_205;
  reg [191:0] _RAND_206;
  reg [191:0] _RAND_207;
  reg [191:0] _RAND_208;
  reg [191:0] _RAND_209;
  reg [191:0] _RAND_210;
  reg [191:0] _RAND_211;
  reg [191:0] _RAND_212;
  reg [191:0] _RAND_213;
  reg [191:0] _RAND_214;
  reg [191:0] _RAND_215;
  reg [191:0] _RAND_216;
  reg [191:0] _RAND_217;
  reg [191:0] _RAND_218;
  reg [191:0] _RAND_219;
  reg [191:0] _RAND_220;
  reg [191:0] _RAND_221;
  reg [191:0] _RAND_222;
  reg [191:0] _RAND_223;
  reg [191:0] _RAND_224;
  reg [191:0] _RAND_225;
  reg [191:0] _RAND_226;
  reg [191:0] _RAND_227;
  reg [191:0] _RAND_228;
  reg [191:0] _RAND_229;
  reg [191:0] _RAND_230;
  reg [191:0] _RAND_231;
  reg [191:0] _RAND_232;
  reg [191:0] _RAND_233;
  reg [191:0] _RAND_234;
  reg [191:0] _RAND_235;
  reg [191:0] _RAND_236;
  reg [191:0] _RAND_237;
  reg [191:0] _RAND_238;
  reg [191:0] _RAND_239;
  reg [191:0] _RAND_240;
  reg [191:0] _RAND_241;
  reg [191:0] _RAND_242;
  reg [191:0] _RAND_243;
  reg [191:0] _RAND_244;
  reg [191:0] _RAND_245;
  reg [191:0] _RAND_246;
  reg [191:0] _RAND_247;
  reg [191:0] _RAND_248;
  reg [191:0] _RAND_249;
  reg [191:0] _RAND_250;
  reg [191:0] _RAND_251;
  reg [191:0] _RAND_252;
  reg [191:0] _RAND_253;
  reg [191:0] _RAND_254;
  reg [191:0] _RAND_255;
  reg [191:0] _RAND_256;
  reg [191:0] _RAND_257;
  reg [191:0] _RAND_258;
  reg [191:0] _RAND_259;
  reg [191:0] _RAND_260;
  reg [191:0] _RAND_261;
  reg [191:0] _RAND_262;
  reg [191:0] _RAND_263;
  reg [191:0] _RAND_264;
  reg [191:0] _RAND_265;
  reg [191:0] _RAND_266;
  reg [191:0] _RAND_267;
  reg [191:0] _RAND_268;
  reg [191:0] _RAND_269;
  reg [191:0] _RAND_270;
  reg [191:0] _RAND_271;
  reg [191:0] _RAND_272;
  reg [191:0] _RAND_273;
  reg [191:0] _RAND_274;
  reg [191:0] _RAND_275;
  reg [191:0] _RAND_276;
  reg [191:0] _RAND_277;
  reg [191:0] _RAND_278;
  reg [191:0] _RAND_279;
  reg [191:0] _RAND_280;
  reg [191:0] _RAND_281;
  reg [191:0] _RAND_282;
  reg [191:0] _RAND_283;
  reg [191:0] _RAND_284;
  reg [191:0] _RAND_285;
  reg [191:0] _RAND_286;
  reg [191:0] _RAND_287;
  reg [191:0] _RAND_288;
  reg [191:0] _RAND_289;
  reg [191:0] _RAND_290;
  reg [191:0] _RAND_291;
  reg [191:0] _RAND_292;
  reg [191:0] _RAND_293;
  reg [191:0] _RAND_294;
  reg [191:0] _RAND_295;
  reg [191:0] _RAND_296;
  reg [191:0] _RAND_297;
  reg [191:0] _RAND_298;
  reg [191:0] _RAND_299;
  reg [191:0] _RAND_300;
  reg [191:0] _RAND_301;
  reg [191:0] _RAND_302;
  reg [191:0] _RAND_303;
  reg [191:0] _RAND_304;
  reg [191:0] _RAND_305;
  reg [191:0] _RAND_306;
  reg [191:0] _RAND_307;
  reg [191:0] _RAND_308;
  reg [191:0] _RAND_309;
  reg [191:0] _RAND_310;
  reg [191:0] _RAND_311;
  reg [191:0] _RAND_312;
  reg [191:0] _RAND_313;
  reg [191:0] _RAND_314;
  reg [191:0] _RAND_315;
  reg [191:0] _RAND_316;
  reg [191:0] _RAND_317;
  reg [191:0] _RAND_318;
  reg [191:0] _RAND_319;
  reg [191:0] _RAND_320;
  reg [191:0] _RAND_321;
  reg [191:0] _RAND_322;
  reg [191:0] _RAND_323;
  reg [191:0] _RAND_324;
  reg [191:0] _RAND_325;
  reg [191:0] _RAND_326;
  reg [191:0] _RAND_327;
  reg [191:0] _RAND_328;
  reg [191:0] _RAND_329;
  reg [191:0] _RAND_330;
  reg [191:0] _RAND_331;
  reg [191:0] _RAND_332;
  reg [191:0] _RAND_333;
  reg [191:0] _RAND_334;
  reg [191:0] _RAND_335;
  reg [191:0] _RAND_336;
  reg [191:0] _RAND_337;
  reg [191:0] _RAND_338;
  reg [191:0] _RAND_339;
  reg [191:0] _RAND_340;
  reg [191:0] _RAND_341;
  reg [191:0] _RAND_342;
  reg [191:0] _RAND_343;
  reg [191:0] _RAND_344;
  reg [191:0] _RAND_345;
  reg [191:0] _RAND_346;
  reg [191:0] _RAND_347;
  reg [191:0] _RAND_348;
  reg [191:0] _RAND_349;
  reg [191:0] _RAND_350;
  reg [191:0] _RAND_351;
  reg [191:0] _RAND_352;
  reg [191:0] _RAND_353;
  reg [191:0] _RAND_354;
  reg [191:0] _RAND_355;
  reg [191:0] _RAND_356;
  reg [191:0] _RAND_357;
  reg [191:0] _RAND_358;
  reg [191:0] _RAND_359;
  reg [191:0] _RAND_360;
  reg [191:0] _RAND_361;
  reg [191:0] _RAND_362;
  reg [191:0] _RAND_363;
  reg [191:0] _RAND_364;
  reg [191:0] _RAND_365;
  reg [191:0] _RAND_366;
  reg [191:0] _RAND_367;
  reg [191:0] _RAND_368;
  reg [191:0] _RAND_369;
  reg [191:0] _RAND_370;
  reg [191:0] _RAND_371;
  reg [191:0] _RAND_372;
  reg [191:0] _RAND_373;
  reg [191:0] _RAND_374;
  reg [191:0] _RAND_375;
  reg [191:0] _RAND_376;
  reg [191:0] _RAND_377;
  reg [191:0] _RAND_378;
  reg [191:0] _RAND_379;
  reg [191:0] _RAND_380;
  reg [191:0] _RAND_381;
  reg [191:0] _RAND_382;
  reg [191:0] _RAND_383;
  reg [191:0] _RAND_384;
  reg [191:0] _RAND_385;
  reg [191:0] _RAND_386;
  reg [191:0] _RAND_387;
  reg [191:0] _RAND_388;
  reg [191:0] _RAND_389;
  reg [191:0] _RAND_390;
  reg [191:0] _RAND_391;
  reg [191:0] _RAND_392;
  reg [191:0] _RAND_393;
  reg [191:0] _RAND_394;
  reg [191:0] _RAND_395;
  reg [191:0] _RAND_396;
  reg [191:0] _RAND_397;
  reg [191:0] _RAND_398;
  reg [191:0] _RAND_399;
  reg [191:0] _RAND_400;
  reg [191:0] _RAND_401;
  reg [191:0] _RAND_402;
  reg [191:0] _RAND_403;
  reg [191:0] _RAND_404;
  reg [191:0] _RAND_405;
  reg [191:0] _RAND_406;
  reg [191:0] _RAND_407;
  reg [191:0] _RAND_408;
  reg [191:0] _RAND_409;
  reg [191:0] _RAND_410;
  reg [191:0] _RAND_411;
  reg [191:0] _RAND_412;
  reg [191:0] _RAND_413;
  reg [191:0] _RAND_414;
  reg [191:0] _RAND_415;
  reg [191:0] _RAND_416;
  reg [191:0] _RAND_417;
  reg [191:0] _RAND_418;
  reg [191:0] _RAND_419;
  reg [191:0] _RAND_420;
  reg [191:0] _RAND_421;
  reg [191:0] _RAND_422;
  reg [191:0] _RAND_423;
  reg [191:0] _RAND_424;
  reg [191:0] _RAND_425;
  reg [191:0] _RAND_426;
  reg [191:0] _RAND_427;
  reg [191:0] _RAND_428;
  reg [191:0] _RAND_429;
  reg [191:0] _RAND_430;
  reg [191:0] _RAND_431;
  reg [191:0] _RAND_432;
  reg [191:0] _RAND_433;
  reg [191:0] _RAND_434;
  reg [191:0] _RAND_435;
  reg [191:0] _RAND_436;
  reg [191:0] _RAND_437;
  reg [191:0] _RAND_438;
  reg [191:0] _RAND_439;
  reg [191:0] _RAND_440;
  reg [191:0] _RAND_441;
  reg [191:0] _RAND_442;
  reg [191:0] _RAND_443;
  reg [191:0] _RAND_444;
  reg [191:0] _RAND_445;
  reg [191:0] _RAND_446;
  reg [191:0] _RAND_447;
  reg [191:0] _RAND_448;
  reg [191:0] _RAND_449;
  reg [191:0] _RAND_450;
  reg [191:0] _RAND_451;
  reg [191:0] _RAND_452;
  reg [191:0] _RAND_453;
  reg [191:0] _RAND_454;
  reg [191:0] _RAND_455;
  reg [191:0] _RAND_456;
  reg [191:0] _RAND_457;
  reg [191:0] _RAND_458;
  reg [191:0] _RAND_459;
  reg [191:0] _RAND_460;
  reg [191:0] _RAND_461;
  reg [191:0] _RAND_462;
  reg [191:0] _RAND_463;
  reg [191:0] _RAND_464;
  reg [191:0] _RAND_465;
  reg [191:0] _RAND_466;
  reg [191:0] _RAND_467;
  reg [191:0] _RAND_468;
  reg [191:0] _RAND_469;
  reg [191:0] _RAND_470;
  reg [191:0] _RAND_471;
  reg [191:0] _RAND_472;
  reg [191:0] _RAND_473;
  reg [191:0] _RAND_474;
  reg [191:0] _RAND_475;
  reg [191:0] _RAND_476;
  reg [191:0] _RAND_477;
  reg [191:0] _RAND_478;
  reg [191:0] _RAND_479;
  reg [191:0] _RAND_480;
  reg [191:0] _RAND_481;
  reg [191:0] _RAND_482;
  reg [191:0] _RAND_483;
  reg [191:0] _RAND_484;
  reg [191:0] _RAND_485;
  reg [191:0] _RAND_486;
  reg [191:0] _RAND_487;
  reg [191:0] _RAND_488;
  reg [191:0] _RAND_489;
  reg [191:0] _RAND_490;
  reg [191:0] _RAND_491;
  reg [191:0] _RAND_492;
  reg [191:0] _RAND_493;
  reg [191:0] _RAND_494;
  reg [191:0] _RAND_495;
  reg [191:0] _RAND_496;
  reg [191:0] _RAND_497;
  reg [191:0] _RAND_498;
  reg [191:0] _RAND_499;
  reg [191:0] _RAND_500;
  reg [191:0] _RAND_501;
  reg [191:0] _RAND_502;
  reg [191:0] _RAND_503;
  reg [191:0] _RAND_504;
  reg [191:0] _RAND_505;
  reg [191:0] _RAND_506;
  reg [191:0] _RAND_507;
  reg [191:0] _RAND_508;
  reg [191:0] _RAND_509;
  reg [191:0] _RAND_510;
  reg [191:0] _RAND_511;
  reg [191:0] _RAND_512;
  reg [191:0] _RAND_513;
  reg [191:0] _RAND_514;
  reg [191:0] _RAND_515;
  reg [191:0] _RAND_516;
  reg [191:0] _RAND_517;
  reg [191:0] _RAND_518;
  reg [191:0] _RAND_519;
  reg [191:0] _RAND_520;
  reg [191:0] _RAND_521;
  reg [191:0] _RAND_522;
  reg [191:0] _RAND_523;
  reg [191:0] _RAND_524;
  reg [191:0] _RAND_525;
  reg [191:0] _RAND_526;
  reg [191:0] _RAND_527;
  reg [191:0] _RAND_528;
  reg [191:0] _RAND_529;
  reg [191:0] _RAND_530;
  reg [191:0] _RAND_531;
  reg [191:0] _RAND_532;
  reg [191:0] _RAND_533;
  reg [191:0] _RAND_534;
  reg [191:0] _RAND_535;
  reg [191:0] _RAND_536;
  reg [191:0] _RAND_537;
  reg [191:0] _RAND_538;
  reg [191:0] _RAND_539;
  reg [191:0] _RAND_540;
  reg [191:0] _RAND_541;
  reg [191:0] _RAND_542;
  reg [191:0] _RAND_543;
  reg [191:0] _RAND_544;
  reg [191:0] _RAND_545;
  reg [191:0] _RAND_546;
  reg [191:0] _RAND_547;
  reg [191:0] _RAND_548;
  reg [191:0] _RAND_549;
  reg [191:0] _RAND_550;
  reg [191:0] _RAND_551;
  reg [191:0] _RAND_552;
  reg [191:0] _RAND_553;
  reg [191:0] _RAND_554;
  reg [191:0] _RAND_555;
  reg [191:0] _RAND_556;
  reg [191:0] _RAND_557;
  reg [191:0] _RAND_558;
  reg [191:0] _RAND_559;
  reg [191:0] _RAND_560;
  reg [191:0] _RAND_561;
  reg [191:0] _RAND_562;
  reg [191:0] _RAND_563;
  reg [191:0] _RAND_564;
  reg [191:0] _RAND_565;
  reg [191:0] _RAND_566;
  reg [191:0] _RAND_567;
  reg [191:0] _RAND_568;
  reg [191:0] _RAND_569;
  reg [191:0] _RAND_570;
  reg [191:0] _RAND_571;
  reg [191:0] _RAND_572;
  reg [191:0] _RAND_573;
  reg [191:0] _RAND_574;
  reg [191:0] _RAND_575;
  reg [191:0] _RAND_576;
  reg [191:0] _RAND_577;
  reg [191:0] _RAND_578;
  reg [191:0] _RAND_579;
  reg [191:0] _RAND_580;
  reg [191:0] _RAND_581;
  reg [191:0] _RAND_582;
  reg [191:0] _RAND_583;
  reg [191:0] _RAND_584;
  reg [191:0] _RAND_585;
  reg [191:0] _RAND_586;
  reg [191:0] _RAND_587;
  reg [191:0] _RAND_588;
  reg [191:0] _RAND_589;
  reg [191:0] _RAND_590;
  reg [191:0] _RAND_591;
  reg [191:0] _RAND_592;
  reg [191:0] _RAND_593;
  reg [191:0] _RAND_594;
  reg [191:0] _RAND_595;
  reg [191:0] _RAND_596;
  reg [191:0] _RAND_597;
  reg [191:0] _RAND_598;
  reg [191:0] _RAND_599;
  reg [191:0] _RAND_600;
  reg [191:0] _RAND_601;
  reg [191:0] _RAND_602;
  reg [191:0] _RAND_603;
  reg [191:0] _RAND_604;
  reg [191:0] _RAND_605;
  reg [191:0] _RAND_606;
  reg [191:0] _RAND_607;
  reg [191:0] _RAND_608;
  reg [191:0] _RAND_609;
  reg [191:0] _RAND_610;
  reg [191:0] _RAND_611;
  reg [191:0] _RAND_612;
  reg [191:0] _RAND_613;
  reg [191:0] _RAND_614;
  reg [191:0] _RAND_615;
  reg [191:0] _RAND_616;
  reg [191:0] _RAND_617;
  reg [191:0] _RAND_618;
  reg [191:0] _RAND_619;
  reg [191:0] _RAND_620;
  reg [191:0] _RAND_621;
  reg [191:0] _RAND_622;
  reg [191:0] _RAND_623;
  reg [191:0] _RAND_624;
  reg [191:0] _RAND_625;
  reg [191:0] _RAND_626;
  reg [191:0] _RAND_627;
  reg [191:0] _RAND_628;
  reg [191:0] _RAND_629;
  reg [191:0] _RAND_630;
  reg [191:0] _RAND_631;
  reg [191:0] _RAND_632;
  reg [191:0] _RAND_633;
  reg [191:0] _RAND_634;
  reg [191:0] _RAND_635;
  reg [191:0] _RAND_636;
  reg [191:0] _RAND_637;
  reg [191:0] _RAND_638;
  reg [191:0] _RAND_639;
  reg [191:0] _RAND_640;
  reg [191:0] _RAND_641;
  reg [191:0] _RAND_642;
  reg [191:0] _RAND_643;
  reg [191:0] _RAND_644;
  reg [191:0] _RAND_645;
  reg [191:0] _RAND_646;
  reg [191:0] _RAND_647;
  reg [191:0] _RAND_648;
  reg [191:0] _RAND_649;
  reg [191:0] _RAND_650;
  reg [191:0] _RAND_651;
  reg [191:0] _RAND_652;
  reg [191:0] _RAND_653;
  reg [191:0] _RAND_654;
  reg [191:0] _RAND_655;
  reg [191:0] _RAND_656;
  reg [191:0] _RAND_657;
  reg [191:0] _RAND_658;
  reg [191:0] _RAND_659;
  reg [191:0] _RAND_660;
  reg [191:0] _RAND_661;
  reg [191:0] _RAND_662;
  reg [191:0] _RAND_663;
  reg [191:0] _RAND_664;
  reg [191:0] _RAND_665;
  reg [191:0] _RAND_666;
  reg [191:0] _RAND_667;
  reg [191:0] _RAND_668;
  reg [191:0] _RAND_669;
  reg [191:0] _RAND_670;
  reg [191:0] _RAND_671;
  reg [191:0] _RAND_672;
  reg [191:0] _RAND_673;
  reg [191:0] _RAND_674;
  reg [191:0] _RAND_675;
  reg [191:0] _RAND_676;
  reg [191:0] _RAND_677;
  reg [191:0] _RAND_678;
  reg [191:0] _RAND_679;
  reg [191:0] _RAND_680;
  reg [191:0] _RAND_681;
  reg [191:0] _RAND_682;
  reg [191:0] _RAND_683;
  reg [191:0] _RAND_684;
  reg [191:0] _RAND_685;
  reg [191:0] _RAND_686;
  reg [191:0] _RAND_687;
  reg [191:0] _RAND_688;
  reg [191:0] _RAND_689;
  reg [191:0] _RAND_690;
  reg [191:0] _RAND_691;
  reg [191:0] _RAND_692;
  reg [191:0] _RAND_693;
  reg [191:0] _RAND_694;
  reg [191:0] _RAND_695;
  reg [191:0] _RAND_696;
  reg [191:0] _RAND_697;
  reg [191:0] _RAND_698;
  reg [191:0] _RAND_699;
  reg [191:0] _RAND_700;
  reg [191:0] _RAND_701;
  reg [191:0] _RAND_702;
  reg [191:0] _RAND_703;
  reg [191:0] _RAND_704;
  reg [191:0] _RAND_705;
  reg [191:0] _RAND_706;
  reg [191:0] _RAND_707;
  reg [191:0] _RAND_708;
  reg [191:0] _RAND_709;
  reg [191:0] _RAND_710;
  reg [191:0] _RAND_711;
  reg [191:0] _RAND_712;
  reg [191:0] _RAND_713;
  reg [191:0] _RAND_714;
  reg [191:0] _RAND_715;
  reg [191:0] _RAND_716;
  reg [191:0] _RAND_717;
  reg [191:0] _RAND_718;
  reg [191:0] _RAND_719;
  reg [191:0] _RAND_720;
  reg [191:0] _RAND_721;
  reg [191:0] _RAND_722;
  reg [191:0] _RAND_723;
  reg [191:0] _RAND_724;
  reg [191:0] _RAND_725;
  reg [191:0] _RAND_726;
  reg [191:0] _RAND_727;
  reg [191:0] _RAND_728;
  reg [191:0] _RAND_729;
  reg [191:0] _RAND_730;
  reg [191:0] _RAND_731;
  reg [191:0] _RAND_732;
  reg [191:0] _RAND_733;
  reg [191:0] _RAND_734;
  reg [191:0] _RAND_735;
  reg [191:0] _RAND_736;
  reg [191:0] _RAND_737;
  reg [191:0] _RAND_738;
  reg [191:0] _RAND_739;
  reg [191:0] _RAND_740;
  reg [191:0] _RAND_741;
  reg [191:0] _RAND_742;
  reg [191:0] _RAND_743;
  reg [191:0] _RAND_744;
  reg [191:0] _RAND_745;
  reg [191:0] _RAND_746;
  reg [191:0] _RAND_747;
  reg [191:0] _RAND_748;
  reg [191:0] _RAND_749;
  reg [191:0] _RAND_750;
  reg [191:0] _RAND_751;
  reg [191:0] _RAND_752;
  reg [191:0] _RAND_753;
  reg [191:0] _RAND_754;
  reg [191:0] _RAND_755;
  reg [191:0] _RAND_756;
  reg [191:0] _RAND_757;
  reg [191:0] _RAND_758;
  reg [191:0] _RAND_759;
  reg [191:0] _RAND_760;
  reg [191:0] _RAND_761;
  reg [191:0] _RAND_762;
  reg [191:0] _RAND_763;
  reg [191:0] _RAND_764;
  reg [191:0] _RAND_765;
  reg [191:0] _RAND_766;
  reg [191:0] _RAND_767;
  reg [191:0] _RAND_768;
  reg [191:0] _RAND_769;
  reg [191:0] _RAND_770;
  reg [191:0] _RAND_771;
  reg [191:0] _RAND_772;
  reg [191:0] _RAND_773;
  reg [191:0] _RAND_774;
  reg [191:0] _RAND_775;
  reg [191:0] _RAND_776;
  reg [191:0] _RAND_777;
  reg [191:0] _RAND_778;
  reg [191:0] _RAND_779;
  reg [191:0] _RAND_780;
  reg [191:0] _RAND_781;
  reg [191:0] _RAND_782;
  reg [191:0] _RAND_783;
  reg [191:0] _RAND_784;
  reg [191:0] _RAND_785;
  reg [191:0] _RAND_786;
  reg [191:0] _RAND_787;
  reg [191:0] _RAND_788;
  reg [191:0] _RAND_789;
  reg [191:0] _RAND_790;
  reg [191:0] _RAND_791;
  reg [191:0] _RAND_792;
  reg [191:0] _RAND_793;
  reg [191:0] _RAND_794;
  reg [191:0] _RAND_795;
  reg [191:0] _RAND_796;
  reg [191:0] _RAND_797;
  reg [191:0] _RAND_798;
  reg [191:0] _RAND_799;
  reg [191:0] _RAND_800;
  reg [191:0] _RAND_801;
  reg [191:0] _RAND_802;
  reg [191:0] _RAND_803;
  reg [191:0] _RAND_804;
  reg [191:0] _RAND_805;
  reg [191:0] _RAND_806;
  reg [191:0] _RAND_807;
  reg [191:0] _RAND_808;
  reg [191:0] _RAND_809;
  reg [191:0] _RAND_810;
  reg [191:0] _RAND_811;
  reg [191:0] _RAND_812;
  reg [191:0] _RAND_813;
  reg [191:0] _RAND_814;
  reg [191:0] _RAND_815;
  reg [191:0] _RAND_816;
  reg [191:0] _RAND_817;
  reg [191:0] _RAND_818;
  reg [191:0] _RAND_819;
  reg [191:0] _RAND_820;
  reg [191:0] _RAND_821;
  reg [191:0] _RAND_822;
  reg [191:0] _RAND_823;
  reg [191:0] _RAND_824;
  reg [191:0] _RAND_825;
  reg [191:0] _RAND_826;
  reg [191:0] _RAND_827;
  reg [191:0] _RAND_828;
  reg [191:0] _RAND_829;
  reg [191:0] _RAND_830;
  reg [191:0] _RAND_831;
  reg [191:0] _RAND_832;
  reg [191:0] _RAND_833;
  reg [191:0] _RAND_834;
  reg [191:0] _RAND_835;
  reg [191:0] _RAND_836;
  reg [191:0] _RAND_837;
  reg [191:0] _RAND_838;
  reg [191:0] _RAND_839;
  reg [191:0] _RAND_840;
  reg [191:0] _RAND_841;
  reg [191:0] _RAND_842;
  reg [191:0] _RAND_843;
  reg [191:0] _RAND_844;
  reg [191:0] _RAND_845;
  reg [191:0] _RAND_846;
  reg [191:0] _RAND_847;
  reg [191:0] _RAND_848;
  reg [191:0] _RAND_849;
  reg [191:0] _RAND_850;
  reg [191:0] _RAND_851;
  reg [191:0] _RAND_852;
  reg [191:0] _RAND_853;
  reg [191:0] _RAND_854;
  reg [191:0] _RAND_855;
  reg [191:0] _RAND_856;
  reg [191:0] _RAND_857;
  reg [191:0] _RAND_858;
  reg [191:0] _RAND_859;
  reg [191:0] _RAND_860;
  reg [191:0] _RAND_861;
  reg [191:0] _RAND_862;
  reg [191:0] _RAND_863;
  reg [191:0] _RAND_864;
  reg [191:0] _RAND_865;
  reg [191:0] _RAND_866;
  reg [191:0] _RAND_867;
  reg [191:0] _RAND_868;
  reg [191:0] _RAND_869;
  reg [191:0] _RAND_870;
  reg [191:0] _RAND_871;
  reg [191:0] _RAND_872;
  reg [191:0] _RAND_873;
  reg [191:0] _RAND_874;
  reg [191:0] _RAND_875;
  reg [191:0] _RAND_876;
  reg [191:0] _RAND_877;
  reg [191:0] _RAND_878;
  reg [191:0] _RAND_879;
  reg [191:0] _RAND_880;
  reg [191:0] _RAND_881;
  reg [191:0] _RAND_882;
  reg [191:0] _RAND_883;
  reg [191:0] _RAND_884;
  reg [191:0] _RAND_885;
  reg [191:0] _RAND_886;
  reg [191:0] _RAND_887;
  reg [191:0] _RAND_888;
  reg [191:0] _RAND_889;
  reg [191:0] _RAND_890;
  reg [191:0] _RAND_891;
  reg [191:0] _RAND_892;
  reg [191:0] _RAND_893;
  reg [191:0] _RAND_894;
  reg [191:0] _RAND_895;
  reg [191:0] _RAND_896;
  reg [191:0] _RAND_897;
  reg [191:0] _RAND_898;
  reg [191:0] _RAND_899;
  reg [191:0] _RAND_900;
  reg [191:0] _RAND_901;
  reg [191:0] _RAND_902;
  reg [191:0] _RAND_903;
  reg [191:0] _RAND_904;
  reg [191:0] _RAND_905;
  reg [191:0] _RAND_906;
  reg [191:0] _RAND_907;
  reg [191:0] _RAND_908;
  reg [191:0] _RAND_909;
  reg [191:0] _RAND_910;
  reg [191:0] _RAND_911;
  reg [191:0] _RAND_912;
  reg [191:0] _RAND_913;
  reg [191:0] _RAND_914;
  reg [191:0] _RAND_915;
  reg [191:0] _RAND_916;
  reg [191:0] _RAND_917;
  reg [191:0] _RAND_918;
  reg [191:0] _RAND_919;
  reg [191:0] _RAND_920;
  reg [191:0] _RAND_921;
  reg [191:0] _RAND_922;
  reg [191:0] _RAND_923;
  reg [191:0] _RAND_924;
  reg [191:0] _RAND_925;
  reg [191:0] _RAND_926;
  reg [191:0] _RAND_927;
  reg [191:0] _RAND_928;
  reg [191:0] _RAND_929;
  reg [191:0] _RAND_930;
  reg [191:0] _RAND_931;
  reg [191:0] _RAND_932;
  reg [191:0] _RAND_933;
  reg [191:0] _RAND_934;
  reg [191:0] _RAND_935;
  reg [191:0] _RAND_936;
  reg [191:0] _RAND_937;
  reg [191:0] _RAND_938;
  reg [191:0] _RAND_939;
  reg [191:0] _RAND_940;
  reg [191:0] _RAND_941;
  reg [191:0] _RAND_942;
  reg [191:0] _RAND_943;
  reg [191:0] _RAND_944;
  reg [191:0] _RAND_945;
  reg [191:0] _RAND_946;
  reg [191:0] _RAND_947;
  reg [191:0] _RAND_948;
  reg [191:0] _RAND_949;
  reg [191:0] _RAND_950;
  reg [191:0] _RAND_951;
  reg [191:0] _RAND_952;
  reg [191:0] _RAND_953;
  reg [191:0] _RAND_954;
  reg [191:0] _RAND_955;
  reg [191:0] _RAND_956;
  reg [191:0] _RAND_957;
  reg [191:0] _RAND_958;
  reg [191:0] _RAND_959;
  reg [191:0] _RAND_960;
  reg [191:0] _RAND_961;
  reg [191:0] _RAND_962;
  reg [191:0] _RAND_963;
  reg [191:0] _RAND_964;
  reg [191:0] _RAND_965;
  reg [191:0] _RAND_966;
  reg [191:0] _RAND_967;
  reg [191:0] _RAND_968;
  reg [191:0] _RAND_969;
  reg [191:0] _RAND_970;
  reg [191:0] _RAND_971;
  reg [191:0] _RAND_972;
  reg [191:0] _RAND_973;
  reg [191:0] _RAND_974;
  reg [191:0] _RAND_975;
  reg [191:0] _RAND_976;
  reg [191:0] _RAND_977;
  reg [191:0] _RAND_978;
  reg [191:0] _RAND_979;
  reg [191:0] _RAND_980;
  reg [191:0] _RAND_981;
  reg [191:0] _RAND_982;
  reg [191:0] _RAND_983;
  reg [191:0] _RAND_984;
  reg [191:0] _RAND_985;
  reg [191:0] _RAND_986;
  reg [191:0] _RAND_987;
  reg [191:0] _RAND_988;
  reg [191:0] _RAND_989;
  reg [191:0] _RAND_990;
  reg [191:0] _RAND_991;
  reg [191:0] _RAND_992;
  reg [191:0] _RAND_993;
  reg [191:0] _RAND_994;
  reg [191:0] _RAND_995;
  reg [191:0] _RAND_996;
  reg [191:0] _RAND_997;
  reg [191:0] _RAND_998;
  reg [191:0] _RAND_999;
  reg [191:0] _RAND_1000;
  reg [191:0] _RAND_1001;
  reg [191:0] _RAND_1002;
  reg [191:0] _RAND_1003;
  reg [191:0] _RAND_1004;
  reg [191:0] _RAND_1005;
  reg [191:0] _RAND_1006;
  reg [191:0] _RAND_1007;
  reg [191:0] _RAND_1008;
  reg [191:0] _RAND_1009;
  reg [191:0] _RAND_1010;
  reg [191:0] _RAND_1011;
  reg [191:0] _RAND_1012;
  reg [191:0] _RAND_1013;
  reg [191:0] _RAND_1014;
  reg [191:0] _RAND_1015;
  reg [191:0] _RAND_1016;
  reg [191:0] _RAND_1017;
  reg [191:0] _RAND_1018;
  reg [191:0] _RAND_1019;
  reg [191:0] _RAND_1020;
  reg [191:0] _RAND_1021;
  reg [191:0] _RAND_1022;
  reg [191:0] _RAND_1023;
  reg [191:0] _RAND_1024;
  reg [191:0] _RAND_1025;
  reg [191:0] _RAND_1026;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[icache.scala 23:67]
  wire  lookup = state == 2'h1; // @[icache.scala 25:66]
  wire  replace = state == 2'h2; // @[icache.scala 26:66]
  wire  refill = state == 2'h3; // @[icache.scala 27:66]
  reg [63:0] reg_rdata; // @[icache.scala 40:26]
  reg  delay; // @[icache.scala 41:25]
  wire [54:0] cpu_tag = io_addr[63:9]; // @[icache.scala 42:24]
  wire [9:0] cpu_index = {io_addr[8:0],1'h0}; // @[Cat.scala 31:58]
  reg [184:0] cache_data_0; // @[icache.scala 47:23]
  reg [184:0] cache_data_1; // @[icache.scala 47:23]
  reg [184:0] cache_data_2; // @[icache.scala 47:23]
  reg [184:0] cache_data_3; // @[icache.scala 47:23]
  reg [184:0] cache_data_4; // @[icache.scala 47:23]
  reg [184:0] cache_data_5; // @[icache.scala 47:23]
  reg [184:0] cache_data_6; // @[icache.scala 47:23]
  reg [184:0] cache_data_7; // @[icache.scala 47:23]
  reg [184:0] cache_data_8; // @[icache.scala 47:23]
  reg [184:0] cache_data_9; // @[icache.scala 47:23]
  reg [184:0] cache_data_10; // @[icache.scala 47:23]
  reg [184:0] cache_data_11; // @[icache.scala 47:23]
  reg [184:0] cache_data_12; // @[icache.scala 47:23]
  reg [184:0] cache_data_13; // @[icache.scala 47:23]
  reg [184:0] cache_data_14; // @[icache.scala 47:23]
  reg [184:0] cache_data_15; // @[icache.scala 47:23]
  reg [184:0] cache_data_16; // @[icache.scala 47:23]
  reg [184:0] cache_data_17; // @[icache.scala 47:23]
  reg [184:0] cache_data_18; // @[icache.scala 47:23]
  reg [184:0] cache_data_19; // @[icache.scala 47:23]
  reg [184:0] cache_data_20; // @[icache.scala 47:23]
  reg [184:0] cache_data_21; // @[icache.scala 47:23]
  reg [184:0] cache_data_22; // @[icache.scala 47:23]
  reg [184:0] cache_data_23; // @[icache.scala 47:23]
  reg [184:0] cache_data_24; // @[icache.scala 47:23]
  reg [184:0] cache_data_25; // @[icache.scala 47:23]
  reg [184:0] cache_data_26; // @[icache.scala 47:23]
  reg [184:0] cache_data_27; // @[icache.scala 47:23]
  reg [184:0] cache_data_28; // @[icache.scala 47:23]
  reg [184:0] cache_data_29; // @[icache.scala 47:23]
  reg [184:0] cache_data_30; // @[icache.scala 47:23]
  reg [184:0] cache_data_31; // @[icache.scala 47:23]
  reg [184:0] cache_data_32; // @[icache.scala 47:23]
  reg [184:0] cache_data_33; // @[icache.scala 47:23]
  reg [184:0] cache_data_34; // @[icache.scala 47:23]
  reg [184:0] cache_data_35; // @[icache.scala 47:23]
  reg [184:0] cache_data_36; // @[icache.scala 47:23]
  reg [184:0] cache_data_37; // @[icache.scala 47:23]
  reg [184:0] cache_data_38; // @[icache.scala 47:23]
  reg [184:0] cache_data_39; // @[icache.scala 47:23]
  reg [184:0] cache_data_40; // @[icache.scala 47:23]
  reg [184:0] cache_data_41; // @[icache.scala 47:23]
  reg [184:0] cache_data_42; // @[icache.scala 47:23]
  reg [184:0] cache_data_43; // @[icache.scala 47:23]
  reg [184:0] cache_data_44; // @[icache.scala 47:23]
  reg [184:0] cache_data_45; // @[icache.scala 47:23]
  reg [184:0] cache_data_46; // @[icache.scala 47:23]
  reg [184:0] cache_data_47; // @[icache.scala 47:23]
  reg [184:0] cache_data_48; // @[icache.scala 47:23]
  reg [184:0] cache_data_49; // @[icache.scala 47:23]
  reg [184:0] cache_data_50; // @[icache.scala 47:23]
  reg [184:0] cache_data_51; // @[icache.scala 47:23]
  reg [184:0] cache_data_52; // @[icache.scala 47:23]
  reg [184:0] cache_data_53; // @[icache.scala 47:23]
  reg [184:0] cache_data_54; // @[icache.scala 47:23]
  reg [184:0] cache_data_55; // @[icache.scala 47:23]
  reg [184:0] cache_data_56; // @[icache.scala 47:23]
  reg [184:0] cache_data_57; // @[icache.scala 47:23]
  reg [184:0] cache_data_58; // @[icache.scala 47:23]
  reg [184:0] cache_data_59; // @[icache.scala 47:23]
  reg [184:0] cache_data_60; // @[icache.scala 47:23]
  reg [184:0] cache_data_61; // @[icache.scala 47:23]
  reg [184:0] cache_data_62; // @[icache.scala 47:23]
  reg [184:0] cache_data_63; // @[icache.scala 47:23]
  reg [184:0] cache_data_64; // @[icache.scala 47:23]
  reg [184:0] cache_data_65; // @[icache.scala 47:23]
  reg [184:0] cache_data_66; // @[icache.scala 47:23]
  reg [184:0] cache_data_67; // @[icache.scala 47:23]
  reg [184:0] cache_data_68; // @[icache.scala 47:23]
  reg [184:0] cache_data_69; // @[icache.scala 47:23]
  reg [184:0] cache_data_70; // @[icache.scala 47:23]
  reg [184:0] cache_data_71; // @[icache.scala 47:23]
  reg [184:0] cache_data_72; // @[icache.scala 47:23]
  reg [184:0] cache_data_73; // @[icache.scala 47:23]
  reg [184:0] cache_data_74; // @[icache.scala 47:23]
  reg [184:0] cache_data_75; // @[icache.scala 47:23]
  reg [184:0] cache_data_76; // @[icache.scala 47:23]
  reg [184:0] cache_data_77; // @[icache.scala 47:23]
  reg [184:0] cache_data_78; // @[icache.scala 47:23]
  reg [184:0] cache_data_79; // @[icache.scala 47:23]
  reg [184:0] cache_data_80; // @[icache.scala 47:23]
  reg [184:0] cache_data_81; // @[icache.scala 47:23]
  reg [184:0] cache_data_82; // @[icache.scala 47:23]
  reg [184:0] cache_data_83; // @[icache.scala 47:23]
  reg [184:0] cache_data_84; // @[icache.scala 47:23]
  reg [184:0] cache_data_85; // @[icache.scala 47:23]
  reg [184:0] cache_data_86; // @[icache.scala 47:23]
  reg [184:0] cache_data_87; // @[icache.scala 47:23]
  reg [184:0] cache_data_88; // @[icache.scala 47:23]
  reg [184:0] cache_data_89; // @[icache.scala 47:23]
  reg [184:0] cache_data_90; // @[icache.scala 47:23]
  reg [184:0] cache_data_91; // @[icache.scala 47:23]
  reg [184:0] cache_data_92; // @[icache.scala 47:23]
  reg [184:0] cache_data_93; // @[icache.scala 47:23]
  reg [184:0] cache_data_94; // @[icache.scala 47:23]
  reg [184:0] cache_data_95; // @[icache.scala 47:23]
  reg [184:0] cache_data_96; // @[icache.scala 47:23]
  reg [184:0] cache_data_97; // @[icache.scala 47:23]
  reg [184:0] cache_data_98; // @[icache.scala 47:23]
  reg [184:0] cache_data_99; // @[icache.scala 47:23]
  reg [184:0] cache_data_100; // @[icache.scala 47:23]
  reg [184:0] cache_data_101; // @[icache.scala 47:23]
  reg [184:0] cache_data_102; // @[icache.scala 47:23]
  reg [184:0] cache_data_103; // @[icache.scala 47:23]
  reg [184:0] cache_data_104; // @[icache.scala 47:23]
  reg [184:0] cache_data_105; // @[icache.scala 47:23]
  reg [184:0] cache_data_106; // @[icache.scala 47:23]
  reg [184:0] cache_data_107; // @[icache.scala 47:23]
  reg [184:0] cache_data_108; // @[icache.scala 47:23]
  reg [184:0] cache_data_109; // @[icache.scala 47:23]
  reg [184:0] cache_data_110; // @[icache.scala 47:23]
  reg [184:0] cache_data_111; // @[icache.scala 47:23]
  reg [184:0] cache_data_112; // @[icache.scala 47:23]
  reg [184:0] cache_data_113; // @[icache.scala 47:23]
  reg [184:0] cache_data_114; // @[icache.scala 47:23]
  reg [184:0] cache_data_115; // @[icache.scala 47:23]
  reg [184:0] cache_data_116; // @[icache.scala 47:23]
  reg [184:0] cache_data_117; // @[icache.scala 47:23]
  reg [184:0] cache_data_118; // @[icache.scala 47:23]
  reg [184:0] cache_data_119; // @[icache.scala 47:23]
  reg [184:0] cache_data_120; // @[icache.scala 47:23]
  reg [184:0] cache_data_121; // @[icache.scala 47:23]
  reg [184:0] cache_data_122; // @[icache.scala 47:23]
  reg [184:0] cache_data_123; // @[icache.scala 47:23]
  reg [184:0] cache_data_124; // @[icache.scala 47:23]
  reg [184:0] cache_data_125; // @[icache.scala 47:23]
  reg [184:0] cache_data_126; // @[icache.scala 47:23]
  reg [184:0] cache_data_127; // @[icache.scala 47:23]
  reg [184:0] cache_data_128; // @[icache.scala 47:23]
  reg [184:0] cache_data_129; // @[icache.scala 47:23]
  reg [184:0] cache_data_130; // @[icache.scala 47:23]
  reg [184:0] cache_data_131; // @[icache.scala 47:23]
  reg [184:0] cache_data_132; // @[icache.scala 47:23]
  reg [184:0] cache_data_133; // @[icache.scala 47:23]
  reg [184:0] cache_data_134; // @[icache.scala 47:23]
  reg [184:0] cache_data_135; // @[icache.scala 47:23]
  reg [184:0] cache_data_136; // @[icache.scala 47:23]
  reg [184:0] cache_data_137; // @[icache.scala 47:23]
  reg [184:0] cache_data_138; // @[icache.scala 47:23]
  reg [184:0] cache_data_139; // @[icache.scala 47:23]
  reg [184:0] cache_data_140; // @[icache.scala 47:23]
  reg [184:0] cache_data_141; // @[icache.scala 47:23]
  reg [184:0] cache_data_142; // @[icache.scala 47:23]
  reg [184:0] cache_data_143; // @[icache.scala 47:23]
  reg [184:0] cache_data_144; // @[icache.scala 47:23]
  reg [184:0] cache_data_145; // @[icache.scala 47:23]
  reg [184:0] cache_data_146; // @[icache.scala 47:23]
  reg [184:0] cache_data_147; // @[icache.scala 47:23]
  reg [184:0] cache_data_148; // @[icache.scala 47:23]
  reg [184:0] cache_data_149; // @[icache.scala 47:23]
  reg [184:0] cache_data_150; // @[icache.scala 47:23]
  reg [184:0] cache_data_151; // @[icache.scala 47:23]
  reg [184:0] cache_data_152; // @[icache.scala 47:23]
  reg [184:0] cache_data_153; // @[icache.scala 47:23]
  reg [184:0] cache_data_154; // @[icache.scala 47:23]
  reg [184:0] cache_data_155; // @[icache.scala 47:23]
  reg [184:0] cache_data_156; // @[icache.scala 47:23]
  reg [184:0] cache_data_157; // @[icache.scala 47:23]
  reg [184:0] cache_data_158; // @[icache.scala 47:23]
  reg [184:0] cache_data_159; // @[icache.scala 47:23]
  reg [184:0] cache_data_160; // @[icache.scala 47:23]
  reg [184:0] cache_data_161; // @[icache.scala 47:23]
  reg [184:0] cache_data_162; // @[icache.scala 47:23]
  reg [184:0] cache_data_163; // @[icache.scala 47:23]
  reg [184:0] cache_data_164; // @[icache.scala 47:23]
  reg [184:0] cache_data_165; // @[icache.scala 47:23]
  reg [184:0] cache_data_166; // @[icache.scala 47:23]
  reg [184:0] cache_data_167; // @[icache.scala 47:23]
  reg [184:0] cache_data_168; // @[icache.scala 47:23]
  reg [184:0] cache_data_169; // @[icache.scala 47:23]
  reg [184:0] cache_data_170; // @[icache.scala 47:23]
  reg [184:0] cache_data_171; // @[icache.scala 47:23]
  reg [184:0] cache_data_172; // @[icache.scala 47:23]
  reg [184:0] cache_data_173; // @[icache.scala 47:23]
  reg [184:0] cache_data_174; // @[icache.scala 47:23]
  reg [184:0] cache_data_175; // @[icache.scala 47:23]
  reg [184:0] cache_data_176; // @[icache.scala 47:23]
  reg [184:0] cache_data_177; // @[icache.scala 47:23]
  reg [184:0] cache_data_178; // @[icache.scala 47:23]
  reg [184:0] cache_data_179; // @[icache.scala 47:23]
  reg [184:0] cache_data_180; // @[icache.scala 47:23]
  reg [184:0] cache_data_181; // @[icache.scala 47:23]
  reg [184:0] cache_data_182; // @[icache.scala 47:23]
  reg [184:0] cache_data_183; // @[icache.scala 47:23]
  reg [184:0] cache_data_184; // @[icache.scala 47:23]
  reg [184:0] cache_data_185; // @[icache.scala 47:23]
  reg [184:0] cache_data_186; // @[icache.scala 47:23]
  reg [184:0] cache_data_187; // @[icache.scala 47:23]
  reg [184:0] cache_data_188; // @[icache.scala 47:23]
  reg [184:0] cache_data_189; // @[icache.scala 47:23]
  reg [184:0] cache_data_190; // @[icache.scala 47:23]
  reg [184:0] cache_data_191; // @[icache.scala 47:23]
  reg [184:0] cache_data_192; // @[icache.scala 47:23]
  reg [184:0] cache_data_193; // @[icache.scala 47:23]
  reg [184:0] cache_data_194; // @[icache.scala 47:23]
  reg [184:0] cache_data_195; // @[icache.scala 47:23]
  reg [184:0] cache_data_196; // @[icache.scala 47:23]
  reg [184:0] cache_data_197; // @[icache.scala 47:23]
  reg [184:0] cache_data_198; // @[icache.scala 47:23]
  reg [184:0] cache_data_199; // @[icache.scala 47:23]
  reg [184:0] cache_data_200; // @[icache.scala 47:23]
  reg [184:0] cache_data_201; // @[icache.scala 47:23]
  reg [184:0] cache_data_202; // @[icache.scala 47:23]
  reg [184:0] cache_data_203; // @[icache.scala 47:23]
  reg [184:0] cache_data_204; // @[icache.scala 47:23]
  reg [184:0] cache_data_205; // @[icache.scala 47:23]
  reg [184:0] cache_data_206; // @[icache.scala 47:23]
  reg [184:0] cache_data_207; // @[icache.scala 47:23]
  reg [184:0] cache_data_208; // @[icache.scala 47:23]
  reg [184:0] cache_data_209; // @[icache.scala 47:23]
  reg [184:0] cache_data_210; // @[icache.scala 47:23]
  reg [184:0] cache_data_211; // @[icache.scala 47:23]
  reg [184:0] cache_data_212; // @[icache.scala 47:23]
  reg [184:0] cache_data_213; // @[icache.scala 47:23]
  reg [184:0] cache_data_214; // @[icache.scala 47:23]
  reg [184:0] cache_data_215; // @[icache.scala 47:23]
  reg [184:0] cache_data_216; // @[icache.scala 47:23]
  reg [184:0] cache_data_217; // @[icache.scala 47:23]
  reg [184:0] cache_data_218; // @[icache.scala 47:23]
  reg [184:0] cache_data_219; // @[icache.scala 47:23]
  reg [184:0] cache_data_220; // @[icache.scala 47:23]
  reg [184:0] cache_data_221; // @[icache.scala 47:23]
  reg [184:0] cache_data_222; // @[icache.scala 47:23]
  reg [184:0] cache_data_223; // @[icache.scala 47:23]
  reg [184:0] cache_data_224; // @[icache.scala 47:23]
  reg [184:0] cache_data_225; // @[icache.scala 47:23]
  reg [184:0] cache_data_226; // @[icache.scala 47:23]
  reg [184:0] cache_data_227; // @[icache.scala 47:23]
  reg [184:0] cache_data_228; // @[icache.scala 47:23]
  reg [184:0] cache_data_229; // @[icache.scala 47:23]
  reg [184:0] cache_data_230; // @[icache.scala 47:23]
  reg [184:0] cache_data_231; // @[icache.scala 47:23]
  reg [184:0] cache_data_232; // @[icache.scala 47:23]
  reg [184:0] cache_data_233; // @[icache.scala 47:23]
  reg [184:0] cache_data_234; // @[icache.scala 47:23]
  reg [184:0] cache_data_235; // @[icache.scala 47:23]
  reg [184:0] cache_data_236; // @[icache.scala 47:23]
  reg [184:0] cache_data_237; // @[icache.scala 47:23]
  reg [184:0] cache_data_238; // @[icache.scala 47:23]
  reg [184:0] cache_data_239; // @[icache.scala 47:23]
  reg [184:0] cache_data_240; // @[icache.scala 47:23]
  reg [184:0] cache_data_241; // @[icache.scala 47:23]
  reg [184:0] cache_data_242; // @[icache.scala 47:23]
  reg [184:0] cache_data_243; // @[icache.scala 47:23]
  reg [184:0] cache_data_244; // @[icache.scala 47:23]
  reg [184:0] cache_data_245; // @[icache.scala 47:23]
  reg [184:0] cache_data_246; // @[icache.scala 47:23]
  reg [184:0] cache_data_247; // @[icache.scala 47:23]
  reg [184:0] cache_data_248; // @[icache.scala 47:23]
  reg [184:0] cache_data_249; // @[icache.scala 47:23]
  reg [184:0] cache_data_250; // @[icache.scala 47:23]
  reg [184:0] cache_data_251; // @[icache.scala 47:23]
  reg [184:0] cache_data_252; // @[icache.scala 47:23]
  reg [184:0] cache_data_253; // @[icache.scala 47:23]
  reg [184:0] cache_data_254; // @[icache.scala 47:23]
  reg [184:0] cache_data_255; // @[icache.scala 47:23]
  reg [184:0] cache_data_256; // @[icache.scala 47:23]
  reg [184:0] cache_data_257; // @[icache.scala 47:23]
  reg [184:0] cache_data_258; // @[icache.scala 47:23]
  reg [184:0] cache_data_259; // @[icache.scala 47:23]
  reg [184:0] cache_data_260; // @[icache.scala 47:23]
  reg [184:0] cache_data_261; // @[icache.scala 47:23]
  reg [184:0] cache_data_262; // @[icache.scala 47:23]
  reg [184:0] cache_data_263; // @[icache.scala 47:23]
  reg [184:0] cache_data_264; // @[icache.scala 47:23]
  reg [184:0] cache_data_265; // @[icache.scala 47:23]
  reg [184:0] cache_data_266; // @[icache.scala 47:23]
  reg [184:0] cache_data_267; // @[icache.scala 47:23]
  reg [184:0] cache_data_268; // @[icache.scala 47:23]
  reg [184:0] cache_data_269; // @[icache.scala 47:23]
  reg [184:0] cache_data_270; // @[icache.scala 47:23]
  reg [184:0] cache_data_271; // @[icache.scala 47:23]
  reg [184:0] cache_data_272; // @[icache.scala 47:23]
  reg [184:0] cache_data_273; // @[icache.scala 47:23]
  reg [184:0] cache_data_274; // @[icache.scala 47:23]
  reg [184:0] cache_data_275; // @[icache.scala 47:23]
  reg [184:0] cache_data_276; // @[icache.scala 47:23]
  reg [184:0] cache_data_277; // @[icache.scala 47:23]
  reg [184:0] cache_data_278; // @[icache.scala 47:23]
  reg [184:0] cache_data_279; // @[icache.scala 47:23]
  reg [184:0] cache_data_280; // @[icache.scala 47:23]
  reg [184:0] cache_data_281; // @[icache.scala 47:23]
  reg [184:0] cache_data_282; // @[icache.scala 47:23]
  reg [184:0] cache_data_283; // @[icache.scala 47:23]
  reg [184:0] cache_data_284; // @[icache.scala 47:23]
  reg [184:0] cache_data_285; // @[icache.scala 47:23]
  reg [184:0] cache_data_286; // @[icache.scala 47:23]
  reg [184:0] cache_data_287; // @[icache.scala 47:23]
  reg [184:0] cache_data_288; // @[icache.scala 47:23]
  reg [184:0] cache_data_289; // @[icache.scala 47:23]
  reg [184:0] cache_data_290; // @[icache.scala 47:23]
  reg [184:0] cache_data_291; // @[icache.scala 47:23]
  reg [184:0] cache_data_292; // @[icache.scala 47:23]
  reg [184:0] cache_data_293; // @[icache.scala 47:23]
  reg [184:0] cache_data_294; // @[icache.scala 47:23]
  reg [184:0] cache_data_295; // @[icache.scala 47:23]
  reg [184:0] cache_data_296; // @[icache.scala 47:23]
  reg [184:0] cache_data_297; // @[icache.scala 47:23]
  reg [184:0] cache_data_298; // @[icache.scala 47:23]
  reg [184:0] cache_data_299; // @[icache.scala 47:23]
  reg [184:0] cache_data_300; // @[icache.scala 47:23]
  reg [184:0] cache_data_301; // @[icache.scala 47:23]
  reg [184:0] cache_data_302; // @[icache.scala 47:23]
  reg [184:0] cache_data_303; // @[icache.scala 47:23]
  reg [184:0] cache_data_304; // @[icache.scala 47:23]
  reg [184:0] cache_data_305; // @[icache.scala 47:23]
  reg [184:0] cache_data_306; // @[icache.scala 47:23]
  reg [184:0] cache_data_307; // @[icache.scala 47:23]
  reg [184:0] cache_data_308; // @[icache.scala 47:23]
  reg [184:0] cache_data_309; // @[icache.scala 47:23]
  reg [184:0] cache_data_310; // @[icache.scala 47:23]
  reg [184:0] cache_data_311; // @[icache.scala 47:23]
  reg [184:0] cache_data_312; // @[icache.scala 47:23]
  reg [184:0] cache_data_313; // @[icache.scala 47:23]
  reg [184:0] cache_data_314; // @[icache.scala 47:23]
  reg [184:0] cache_data_315; // @[icache.scala 47:23]
  reg [184:0] cache_data_316; // @[icache.scala 47:23]
  reg [184:0] cache_data_317; // @[icache.scala 47:23]
  reg [184:0] cache_data_318; // @[icache.scala 47:23]
  reg [184:0] cache_data_319; // @[icache.scala 47:23]
  reg [184:0] cache_data_320; // @[icache.scala 47:23]
  reg [184:0] cache_data_321; // @[icache.scala 47:23]
  reg [184:0] cache_data_322; // @[icache.scala 47:23]
  reg [184:0] cache_data_323; // @[icache.scala 47:23]
  reg [184:0] cache_data_324; // @[icache.scala 47:23]
  reg [184:0] cache_data_325; // @[icache.scala 47:23]
  reg [184:0] cache_data_326; // @[icache.scala 47:23]
  reg [184:0] cache_data_327; // @[icache.scala 47:23]
  reg [184:0] cache_data_328; // @[icache.scala 47:23]
  reg [184:0] cache_data_329; // @[icache.scala 47:23]
  reg [184:0] cache_data_330; // @[icache.scala 47:23]
  reg [184:0] cache_data_331; // @[icache.scala 47:23]
  reg [184:0] cache_data_332; // @[icache.scala 47:23]
  reg [184:0] cache_data_333; // @[icache.scala 47:23]
  reg [184:0] cache_data_334; // @[icache.scala 47:23]
  reg [184:0] cache_data_335; // @[icache.scala 47:23]
  reg [184:0] cache_data_336; // @[icache.scala 47:23]
  reg [184:0] cache_data_337; // @[icache.scala 47:23]
  reg [184:0] cache_data_338; // @[icache.scala 47:23]
  reg [184:0] cache_data_339; // @[icache.scala 47:23]
  reg [184:0] cache_data_340; // @[icache.scala 47:23]
  reg [184:0] cache_data_341; // @[icache.scala 47:23]
  reg [184:0] cache_data_342; // @[icache.scala 47:23]
  reg [184:0] cache_data_343; // @[icache.scala 47:23]
  reg [184:0] cache_data_344; // @[icache.scala 47:23]
  reg [184:0] cache_data_345; // @[icache.scala 47:23]
  reg [184:0] cache_data_346; // @[icache.scala 47:23]
  reg [184:0] cache_data_347; // @[icache.scala 47:23]
  reg [184:0] cache_data_348; // @[icache.scala 47:23]
  reg [184:0] cache_data_349; // @[icache.scala 47:23]
  reg [184:0] cache_data_350; // @[icache.scala 47:23]
  reg [184:0] cache_data_351; // @[icache.scala 47:23]
  reg [184:0] cache_data_352; // @[icache.scala 47:23]
  reg [184:0] cache_data_353; // @[icache.scala 47:23]
  reg [184:0] cache_data_354; // @[icache.scala 47:23]
  reg [184:0] cache_data_355; // @[icache.scala 47:23]
  reg [184:0] cache_data_356; // @[icache.scala 47:23]
  reg [184:0] cache_data_357; // @[icache.scala 47:23]
  reg [184:0] cache_data_358; // @[icache.scala 47:23]
  reg [184:0] cache_data_359; // @[icache.scala 47:23]
  reg [184:0] cache_data_360; // @[icache.scala 47:23]
  reg [184:0] cache_data_361; // @[icache.scala 47:23]
  reg [184:0] cache_data_362; // @[icache.scala 47:23]
  reg [184:0] cache_data_363; // @[icache.scala 47:23]
  reg [184:0] cache_data_364; // @[icache.scala 47:23]
  reg [184:0] cache_data_365; // @[icache.scala 47:23]
  reg [184:0] cache_data_366; // @[icache.scala 47:23]
  reg [184:0] cache_data_367; // @[icache.scala 47:23]
  reg [184:0] cache_data_368; // @[icache.scala 47:23]
  reg [184:0] cache_data_369; // @[icache.scala 47:23]
  reg [184:0] cache_data_370; // @[icache.scala 47:23]
  reg [184:0] cache_data_371; // @[icache.scala 47:23]
  reg [184:0] cache_data_372; // @[icache.scala 47:23]
  reg [184:0] cache_data_373; // @[icache.scala 47:23]
  reg [184:0] cache_data_374; // @[icache.scala 47:23]
  reg [184:0] cache_data_375; // @[icache.scala 47:23]
  reg [184:0] cache_data_376; // @[icache.scala 47:23]
  reg [184:0] cache_data_377; // @[icache.scala 47:23]
  reg [184:0] cache_data_378; // @[icache.scala 47:23]
  reg [184:0] cache_data_379; // @[icache.scala 47:23]
  reg [184:0] cache_data_380; // @[icache.scala 47:23]
  reg [184:0] cache_data_381; // @[icache.scala 47:23]
  reg [184:0] cache_data_382; // @[icache.scala 47:23]
  reg [184:0] cache_data_383; // @[icache.scala 47:23]
  reg [184:0] cache_data_384; // @[icache.scala 47:23]
  reg [184:0] cache_data_385; // @[icache.scala 47:23]
  reg [184:0] cache_data_386; // @[icache.scala 47:23]
  reg [184:0] cache_data_387; // @[icache.scala 47:23]
  reg [184:0] cache_data_388; // @[icache.scala 47:23]
  reg [184:0] cache_data_389; // @[icache.scala 47:23]
  reg [184:0] cache_data_390; // @[icache.scala 47:23]
  reg [184:0] cache_data_391; // @[icache.scala 47:23]
  reg [184:0] cache_data_392; // @[icache.scala 47:23]
  reg [184:0] cache_data_393; // @[icache.scala 47:23]
  reg [184:0] cache_data_394; // @[icache.scala 47:23]
  reg [184:0] cache_data_395; // @[icache.scala 47:23]
  reg [184:0] cache_data_396; // @[icache.scala 47:23]
  reg [184:0] cache_data_397; // @[icache.scala 47:23]
  reg [184:0] cache_data_398; // @[icache.scala 47:23]
  reg [184:0] cache_data_399; // @[icache.scala 47:23]
  reg [184:0] cache_data_400; // @[icache.scala 47:23]
  reg [184:0] cache_data_401; // @[icache.scala 47:23]
  reg [184:0] cache_data_402; // @[icache.scala 47:23]
  reg [184:0] cache_data_403; // @[icache.scala 47:23]
  reg [184:0] cache_data_404; // @[icache.scala 47:23]
  reg [184:0] cache_data_405; // @[icache.scala 47:23]
  reg [184:0] cache_data_406; // @[icache.scala 47:23]
  reg [184:0] cache_data_407; // @[icache.scala 47:23]
  reg [184:0] cache_data_408; // @[icache.scala 47:23]
  reg [184:0] cache_data_409; // @[icache.scala 47:23]
  reg [184:0] cache_data_410; // @[icache.scala 47:23]
  reg [184:0] cache_data_411; // @[icache.scala 47:23]
  reg [184:0] cache_data_412; // @[icache.scala 47:23]
  reg [184:0] cache_data_413; // @[icache.scala 47:23]
  reg [184:0] cache_data_414; // @[icache.scala 47:23]
  reg [184:0] cache_data_415; // @[icache.scala 47:23]
  reg [184:0] cache_data_416; // @[icache.scala 47:23]
  reg [184:0] cache_data_417; // @[icache.scala 47:23]
  reg [184:0] cache_data_418; // @[icache.scala 47:23]
  reg [184:0] cache_data_419; // @[icache.scala 47:23]
  reg [184:0] cache_data_420; // @[icache.scala 47:23]
  reg [184:0] cache_data_421; // @[icache.scala 47:23]
  reg [184:0] cache_data_422; // @[icache.scala 47:23]
  reg [184:0] cache_data_423; // @[icache.scala 47:23]
  reg [184:0] cache_data_424; // @[icache.scala 47:23]
  reg [184:0] cache_data_425; // @[icache.scala 47:23]
  reg [184:0] cache_data_426; // @[icache.scala 47:23]
  reg [184:0] cache_data_427; // @[icache.scala 47:23]
  reg [184:0] cache_data_428; // @[icache.scala 47:23]
  reg [184:0] cache_data_429; // @[icache.scala 47:23]
  reg [184:0] cache_data_430; // @[icache.scala 47:23]
  reg [184:0] cache_data_431; // @[icache.scala 47:23]
  reg [184:0] cache_data_432; // @[icache.scala 47:23]
  reg [184:0] cache_data_433; // @[icache.scala 47:23]
  reg [184:0] cache_data_434; // @[icache.scala 47:23]
  reg [184:0] cache_data_435; // @[icache.scala 47:23]
  reg [184:0] cache_data_436; // @[icache.scala 47:23]
  reg [184:0] cache_data_437; // @[icache.scala 47:23]
  reg [184:0] cache_data_438; // @[icache.scala 47:23]
  reg [184:0] cache_data_439; // @[icache.scala 47:23]
  reg [184:0] cache_data_440; // @[icache.scala 47:23]
  reg [184:0] cache_data_441; // @[icache.scala 47:23]
  reg [184:0] cache_data_442; // @[icache.scala 47:23]
  reg [184:0] cache_data_443; // @[icache.scala 47:23]
  reg [184:0] cache_data_444; // @[icache.scala 47:23]
  reg [184:0] cache_data_445; // @[icache.scala 47:23]
  reg [184:0] cache_data_446; // @[icache.scala 47:23]
  reg [184:0] cache_data_447; // @[icache.scala 47:23]
  reg [184:0] cache_data_448; // @[icache.scala 47:23]
  reg [184:0] cache_data_449; // @[icache.scala 47:23]
  reg [184:0] cache_data_450; // @[icache.scala 47:23]
  reg [184:0] cache_data_451; // @[icache.scala 47:23]
  reg [184:0] cache_data_452; // @[icache.scala 47:23]
  reg [184:0] cache_data_453; // @[icache.scala 47:23]
  reg [184:0] cache_data_454; // @[icache.scala 47:23]
  reg [184:0] cache_data_455; // @[icache.scala 47:23]
  reg [184:0] cache_data_456; // @[icache.scala 47:23]
  reg [184:0] cache_data_457; // @[icache.scala 47:23]
  reg [184:0] cache_data_458; // @[icache.scala 47:23]
  reg [184:0] cache_data_459; // @[icache.scala 47:23]
  reg [184:0] cache_data_460; // @[icache.scala 47:23]
  reg [184:0] cache_data_461; // @[icache.scala 47:23]
  reg [184:0] cache_data_462; // @[icache.scala 47:23]
  reg [184:0] cache_data_463; // @[icache.scala 47:23]
  reg [184:0] cache_data_464; // @[icache.scala 47:23]
  reg [184:0] cache_data_465; // @[icache.scala 47:23]
  reg [184:0] cache_data_466; // @[icache.scala 47:23]
  reg [184:0] cache_data_467; // @[icache.scala 47:23]
  reg [184:0] cache_data_468; // @[icache.scala 47:23]
  reg [184:0] cache_data_469; // @[icache.scala 47:23]
  reg [184:0] cache_data_470; // @[icache.scala 47:23]
  reg [184:0] cache_data_471; // @[icache.scala 47:23]
  reg [184:0] cache_data_472; // @[icache.scala 47:23]
  reg [184:0] cache_data_473; // @[icache.scala 47:23]
  reg [184:0] cache_data_474; // @[icache.scala 47:23]
  reg [184:0] cache_data_475; // @[icache.scala 47:23]
  reg [184:0] cache_data_476; // @[icache.scala 47:23]
  reg [184:0] cache_data_477; // @[icache.scala 47:23]
  reg [184:0] cache_data_478; // @[icache.scala 47:23]
  reg [184:0] cache_data_479; // @[icache.scala 47:23]
  reg [184:0] cache_data_480; // @[icache.scala 47:23]
  reg [184:0] cache_data_481; // @[icache.scala 47:23]
  reg [184:0] cache_data_482; // @[icache.scala 47:23]
  reg [184:0] cache_data_483; // @[icache.scala 47:23]
  reg [184:0] cache_data_484; // @[icache.scala 47:23]
  reg [184:0] cache_data_485; // @[icache.scala 47:23]
  reg [184:0] cache_data_486; // @[icache.scala 47:23]
  reg [184:0] cache_data_487; // @[icache.scala 47:23]
  reg [184:0] cache_data_488; // @[icache.scala 47:23]
  reg [184:0] cache_data_489; // @[icache.scala 47:23]
  reg [184:0] cache_data_490; // @[icache.scala 47:23]
  reg [184:0] cache_data_491; // @[icache.scala 47:23]
  reg [184:0] cache_data_492; // @[icache.scala 47:23]
  reg [184:0] cache_data_493; // @[icache.scala 47:23]
  reg [184:0] cache_data_494; // @[icache.scala 47:23]
  reg [184:0] cache_data_495; // @[icache.scala 47:23]
  reg [184:0] cache_data_496; // @[icache.scala 47:23]
  reg [184:0] cache_data_497; // @[icache.scala 47:23]
  reg [184:0] cache_data_498; // @[icache.scala 47:23]
  reg [184:0] cache_data_499; // @[icache.scala 47:23]
  reg [184:0] cache_data_500; // @[icache.scala 47:23]
  reg [184:0] cache_data_501; // @[icache.scala 47:23]
  reg [184:0] cache_data_502; // @[icache.scala 47:23]
  reg [184:0] cache_data_503; // @[icache.scala 47:23]
  reg [184:0] cache_data_504; // @[icache.scala 47:23]
  reg [184:0] cache_data_505; // @[icache.scala 47:23]
  reg [184:0] cache_data_506; // @[icache.scala 47:23]
  reg [184:0] cache_data_507; // @[icache.scala 47:23]
  reg [184:0] cache_data_508; // @[icache.scala 47:23]
  reg [184:0] cache_data_509; // @[icache.scala 47:23]
  reg [184:0] cache_data_510; // @[icache.scala 47:23]
  reg [184:0] cache_data_511; // @[icache.scala 47:23]
  reg [184:0] cache_data_512; // @[icache.scala 47:23]
  reg [184:0] cache_data_513; // @[icache.scala 47:23]
  reg [184:0] cache_data_514; // @[icache.scala 47:23]
  reg [184:0] cache_data_515; // @[icache.scala 47:23]
  reg [184:0] cache_data_516; // @[icache.scala 47:23]
  reg [184:0] cache_data_517; // @[icache.scala 47:23]
  reg [184:0] cache_data_518; // @[icache.scala 47:23]
  reg [184:0] cache_data_519; // @[icache.scala 47:23]
  reg [184:0] cache_data_520; // @[icache.scala 47:23]
  reg [184:0] cache_data_521; // @[icache.scala 47:23]
  reg [184:0] cache_data_522; // @[icache.scala 47:23]
  reg [184:0] cache_data_523; // @[icache.scala 47:23]
  reg [184:0] cache_data_524; // @[icache.scala 47:23]
  reg [184:0] cache_data_525; // @[icache.scala 47:23]
  reg [184:0] cache_data_526; // @[icache.scala 47:23]
  reg [184:0] cache_data_527; // @[icache.scala 47:23]
  reg [184:0] cache_data_528; // @[icache.scala 47:23]
  reg [184:0] cache_data_529; // @[icache.scala 47:23]
  reg [184:0] cache_data_530; // @[icache.scala 47:23]
  reg [184:0] cache_data_531; // @[icache.scala 47:23]
  reg [184:0] cache_data_532; // @[icache.scala 47:23]
  reg [184:0] cache_data_533; // @[icache.scala 47:23]
  reg [184:0] cache_data_534; // @[icache.scala 47:23]
  reg [184:0] cache_data_535; // @[icache.scala 47:23]
  reg [184:0] cache_data_536; // @[icache.scala 47:23]
  reg [184:0] cache_data_537; // @[icache.scala 47:23]
  reg [184:0] cache_data_538; // @[icache.scala 47:23]
  reg [184:0] cache_data_539; // @[icache.scala 47:23]
  reg [184:0] cache_data_540; // @[icache.scala 47:23]
  reg [184:0] cache_data_541; // @[icache.scala 47:23]
  reg [184:0] cache_data_542; // @[icache.scala 47:23]
  reg [184:0] cache_data_543; // @[icache.scala 47:23]
  reg [184:0] cache_data_544; // @[icache.scala 47:23]
  reg [184:0] cache_data_545; // @[icache.scala 47:23]
  reg [184:0] cache_data_546; // @[icache.scala 47:23]
  reg [184:0] cache_data_547; // @[icache.scala 47:23]
  reg [184:0] cache_data_548; // @[icache.scala 47:23]
  reg [184:0] cache_data_549; // @[icache.scala 47:23]
  reg [184:0] cache_data_550; // @[icache.scala 47:23]
  reg [184:0] cache_data_551; // @[icache.scala 47:23]
  reg [184:0] cache_data_552; // @[icache.scala 47:23]
  reg [184:0] cache_data_553; // @[icache.scala 47:23]
  reg [184:0] cache_data_554; // @[icache.scala 47:23]
  reg [184:0] cache_data_555; // @[icache.scala 47:23]
  reg [184:0] cache_data_556; // @[icache.scala 47:23]
  reg [184:0] cache_data_557; // @[icache.scala 47:23]
  reg [184:0] cache_data_558; // @[icache.scala 47:23]
  reg [184:0] cache_data_559; // @[icache.scala 47:23]
  reg [184:0] cache_data_560; // @[icache.scala 47:23]
  reg [184:0] cache_data_561; // @[icache.scala 47:23]
  reg [184:0] cache_data_562; // @[icache.scala 47:23]
  reg [184:0] cache_data_563; // @[icache.scala 47:23]
  reg [184:0] cache_data_564; // @[icache.scala 47:23]
  reg [184:0] cache_data_565; // @[icache.scala 47:23]
  reg [184:0] cache_data_566; // @[icache.scala 47:23]
  reg [184:0] cache_data_567; // @[icache.scala 47:23]
  reg [184:0] cache_data_568; // @[icache.scala 47:23]
  reg [184:0] cache_data_569; // @[icache.scala 47:23]
  reg [184:0] cache_data_570; // @[icache.scala 47:23]
  reg [184:0] cache_data_571; // @[icache.scala 47:23]
  reg [184:0] cache_data_572; // @[icache.scala 47:23]
  reg [184:0] cache_data_573; // @[icache.scala 47:23]
  reg [184:0] cache_data_574; // @[icache.scala 47:23]
  reg [184:0] cache_data_575; // @[icache.scala 47:23]
  reg [184:0] cache_data_576; // @[icache.scala 47:23]
  reg [184:0] cache_data_577; // @[icache.scala 47:23]
  reg [184:0] cache_data_578; // @[icache.scala 47:23]
  reg [184:0] cache_data_579; // @[icache.scala 47:23]
  reg [184:0] cache_data_580; // @[icache.scala 47:23]
  reg [184:0] cache_data_581; // @[icache.scala 47:23]
  reg [184:0] cache_data_582; // @[icache.scala 47:23]
  reg [184:0] cache_data_583; // @[icache.scala 47:23]
  reg [184:0] cache_data_584; // @[icache.scala 47:23]
  reg [184:0] cache_data_585; // @[icache.scala 47:23]
  reg [184:0] cache_data_586; // @[icache.scala 47:23]
  reg [184:0] cache_data_587; // @[icache.scala 47:23]
  reg [184:0] cache_data_588; // @[icache.scala 47:23]
  reg [184:0] cache_data_589; // @[icache.scala 47:23]
  reg [184:0] cache_data_590; // @[icache.scala 47:23]
  reg [184:0] cache_data_591; // @[icache.scala 47:23]
  reg [184:0] cache_data_592; // @[icache.scala 47:23]
  reg [184:0] cache_data_593; // @[icache.scala 47:23]
  reg [184:0] cache_data_594; // @[icache.scala 47:23]
  reg [184:0] cache_data_595; // @[icache.scala 47:23]
  reg [184:0] cache_data_596; // @[icache.scala 47:23]
  reg [184:0] cache_data_597; // @[icache.scala 47:23]
  reg [184:0] cache_data_598; // @[icache.scala 47:23]
  reg [184:0] cache_data_599; // @[icache.scala 47:23]
  reg [184:0] cache_data_600; // @[icache.scala 47:23]
  reg [184:0] cache_data_601; // @[icache.scala 47:23]
  reg [184:0] cache_data_602; // @[icache.scala 47:23]
  reg [184:0] cache_data_603; // @[icache.scala 47:23]
  reg [184:0] cache_data_604; // @[icache.scala 47:23]
  reg [184:0] cache_data_605; // @[icache.scala 47:23]
  reg [184:0] cache_data_606; // @[icache.scala 47:23]
  reg [184:0] cache_data_607; // @[icache.scala 47:23]
  reg [184:0] cache_data_608; // @[icache.scala 47:23]
  reg [184:0] cache_data_609; // @[icache.scala 47:23]
  reg [184:0] cache_data_610; // @[icache.scala 47:23]
  reg [184:0] cache_data_611; // @[icache.scala 47:23]
  reg [184:0] cache_data_612; // @[icache.scala 47:23]
  reg [184:0] cache_data_613; // @[icache.scala 47:23]
  reg [184:0] cache_data_614; // @[icache.scala 47:23]
  reg [184:0] cache_data_615; // @[icache.scala 47:23]
  reg [184:0] cache_data_616; // @[icache.scala 47:23]
  reg [184:0] cache_data_617; // @[icache.scala 47:23]
  reg [184:0] cache_data_618; // @[icache.scala 47:23]
  reg [184:0] cache_data_619; // @[icache.scala 47:23]
  reg [184:0] cache_data_620; // @[icache.scala 47:23]
  reg [184:0] cache_data_621; // @[icache.scala 47:23]
  reg [184:0] cache_data_622; // @[icache.scala 47:23]
  reg [184:0] cache_data_623; // @[icache.scala 47:23]
  reg [184:0] cache_data_624; // @[icache.scala 47:23]
  reg [184:0] cache_data_625; // @[icache.scala 47:23]
  reg [184:0] cache_data_626; // @[icache.scala 47:23]
  reg [184:0] cache_data_627; // @[icache.scala 47:23]
  reg [184:0] cache_data_628; // @[icache.scala 47:23]
  reg [184:0] cache_data_629; // @[icache.scala 47:23]
  reg [184:0] cache_data_630; // @[icache.scala 47:23]
  reg [184:0] cache_data_631; // @[icache.scala 47:23]
  reg [184:0] cache_data_632; // @[icache.scala 47:23]
  reg [184:0] cache_data_633; // @[icache.scala 47:23]
  reg [184:0] cache_data_634; // @[icache.scala 47:23]
  reg [184:0] cache_data_635; // @[icache.scala 47:23]
  reg [184:0] cache_data_636; // @[icache.scala 47:23]
  reg [184:0] cache_data_637; // @[icache.scala 47:23]
  reg [184:0] cache_data_638; // @[icache.scala 47:23]
  reg [184:0] cache_data_639; // @[icache.scala 47:23]
  reg [184:0] cache_data_640; // @[icache.scala 47:23]
  reg [184:0] cache_data_641; // @[icache.scala 47:23]
  reg [184:0] cache_data_642; // @[icache.scala 47:23]
  reg [184:0] cache_data_643; // @[icache.scala 47:23]
  reg [184:0] cache_data_644; // @[icache.scala 47:23]
  reg [184:0] cache_data_645; // @[icache.scala 47:23]
  reg [184:0] cache_data_646; // @[icache.scala 47:23]
  reg [184:0] cache_data_647; // @[icache.scala 47:23]
  reg [184:0] cache_data_648; // @[icache.scala 47:23]
  reg [184:0] cache_data_649; // @[icache.scala 47:23]
  reg [184:0] cache_data_650; // @[icache.scala 47:23]
  reg [184:0] cache_data_651; // @[icache.scala 47:23]
  reg [184:0] cache_data_652; // @[icache.scala 47:23]
  reg [184:0] cache_data_653; // @[icache.scala 47:23]
  reg [184:0] cache_data_654; // @[icache.scala 47:23]
  reg [184:0] cache_data_655; // @[icache.scala 47:23]
  reg [184:0] cache_data_656; // @[icache.scala 47:23]
  reg [184:0] cache_data_657; // @[icache.scala 47:23]
  reg [184:0] cache_data_658; // @[icache.scala 47:23]
  reg [184:0] cache_data_659; // @[icache.scala 47:23]
  reg [184:0] cache_data_660; // @[icache.scala 47:23]
  reg [184:0] cache_data_661; // @[icache.scala 47:23]
  reg [184:0] cache_data_662; // @[icache.scala 47:23]
  reg [184:0] cache_data_663; // @[icache.scala 47:23]
  reg [184:0] cache_data_664; // @[icache.scala 47:23]
  reg [184:0] cache_data_665; // @[icache.scala 47:23]
  reg [184:0] cache_data_666; // @[icache.scala 47:23]
  reg [184:0] cache_data_667; // @[icache.scala 47:23]
  reg [184:0] cache_data_668; // @[icache.scala 47:23]
  reg [184:0] cache_data_669; // @[icache.scala 47:23]
  reg [184:0] cache_data_670; // @[icache.scala 47:23]
  reg [184:0] cache_data_671; // @[icache.scala 47:23]
  reg [184:0] cache_data_672; // @[icache.scala 47:23]
  reg [184:0] cache_data_673; // @[icache.scala 47:23]
  reg [184:0] cache_data_674; // @[icache.scala 47:23]
  reg [184:0] cache_data_675; // @[icache.scala 47:23]
  reg [184:0] cache_data_676; // @[icache.scala 47:23]
  reg [184:0] cache_data_677; // @[icache.scala 47:23]
  reg [184:0] cache_data_678; // @[icache.scala 47:23]
  reg [184:0] cache_data_679; // @[icache.scala 47:23]
  reg [184:0] cache_data_680; // @[icache.scala 47:23]
  reg [184:0] cache_data_681; // @[icache.scala 47:23]
  reg [184:0] cache_data_682; // @[icache.scala 47:23]
  reg [184:0] cache_data_683; // @[icache.scala 47:23]
  reg [184:0] cache_data_684; // @[icache.scala 47:23]
  reg [184:0] cache_data_685; // @[icache.scala 47:23]
  reg [184:0] cache_data_686; // @[icache.scala 47:23]
  reg [184:0] cache_data_687; // @[icache.scala 47:23]
  reg [184:0] cache_data_688; // @[icache.scala 47:23]
  reg [184:0] cache_data_689; // @[icache.scala 47:23]
  reg [184:0] cache_data_690; // @[icache.scala 47:23]
  reg [184:0] cache_data_691; // @[icache.scala 47:23]
  reg [184:0] cache_data_692; // @[icache.scala 47:23]
  reg [184:0] cache_data_693; // @[icache.scala 47:23]
  reg [184:0] cache_data_694; // @[icache.scala 47:23]
  reg [184:0] cache_data_695; // @[icache.scala 47:23]
  reg [184:0] cache_data_696; // @[icache.scala 47:23]
  reg [184:0] cache_data_697; // @[icache.scala 47:23]
  reg [184:0] cache_data_698; // @[icache.scala 47:23]
  reg [184:0] cache_data_699; // @[icache.scala 47:23]
  reg [184:0] cache_data_700; // @[icache.scala 47:23]
  reg [184:0] cache_data_701; // @[icache.scala 47:23]
  reg [184:0] cache_data_702; // @[icache.scala 47:23]
  reg [184:0] cache_data_703; // @[icache.scala 47:23]
  reg [184:0] cache_data_704; // @[icache.scala 47:23]
  reg [184:0] cache_data_705; // @[icache.scala 47:23]
  reg [184:0] cache_data_706; // @[icache.scala 47:23]
  reg [184:0] cache_data_707; // @[icache.scala 47:23]
  reg [184:0] cache_data_708; // @[icache.scala 47:23]
  reg [184:0] cache_data_709; // @[icache.scala 47:23]
  reg [184:0] cache_data_710; // @[icache.scala 47:23]
  reg [184:0] cache_data_711; // @[icache.scala 47:23]
  reg [184:0] cache_data_712; // @[icache.scala 47:23]
  reg [184:0] cache_data_713; // @[icache.scala 47:23]
  reg [184:0] cache_data_714; // @[icache.scala 47:23]
  reg [184:0] cache_data_715; // @[icache.scala 47:23]
  reg [184:0] cache_data_716; // @[icache.scala 47:23]
  reg [184:0] cache_data_717; // @[icache.scala 47:23]
  reg [184:0] cache_data_718; // @[icache.scala 47:23]
  reg [184:0] cache_data_719; // @[icache.scala 47:23]
  reg [184:0] cache_data_720; // @[icache.scala 47:23]
  reg [184:0] cache_data_721; // @[icache.scala 47:23]
  reg [184:0] cache_data_722; // @[icache.scala 47:23]
  reg [184:0] cache_data_723; // @[icache.scala 47:23]
  reg [184:0] cache_data_724; // @[icache.scala 47:23]
  reg [184:0] cache_data_725; // @[icache.scala 47:23]
  reg [184:0] cache_data_726; // @[icache.scala 47:23]
  reg [184:0] cache_data_727; // @[icache.scala 47:23]
  reg [184:0] cache_data_728; // @[icache.scala 47:23]
  reg [184:0] cache_data_729; // @[icache.scala 47:23]
  reg [184:0] cache_data_730; // @[icache.scala 47:23]
  reg [184:0] cache_data_731; // @[icache.scala 47:23]
  reg [184:0] cache_data_732; // @[icache.scala 47:23]
  reg [184:0] cache_data_733; // @[icache.scala 47:23]
  reg [184:0] cache_data_734; // @[icache.scala 47:23]
  reg [184:0] cache_data_735; // @[icache.scala 47:23]
  reg [184:0] cache_data_736; // @[icache.scala 47:23]
  reg [184:0] cache_data_737; // @[icache.scala 47:23]
  reg [184:0] cache_data_738; // @[icache.scala 47:23]
  reg [184:0] cache_data_739; // @[icache.scala 47:23]
  reg [184:0] cache_data_740; // @[icache.scala 47:23]
  reg [184:0] cache_data_741; // @[icache.scala 47:23]
  reg [184:0] cache_data_742; // @[icache.scala 47:23]
  reg [184:0] cache_data_743; // @[icache.scala 47:23]
  reg [184:0] cache_data_744; // @[icache.scala 47:23]
  reg [184:0] cache_data_745; // @[icache.scala 47:23]
  reg [184:0] cache_data_746; // @[icache.scala 47:23]
  reg [184:0] cache_data_747; // @[icache.scala 47:23]
  reg [184:0] cache_data_748; // @[icache.scala 47:23]
  reg [184:0] cache_data_749; // @[icache.scala 47:23]
  reg [184:0] cache_data_750; // @[icache.scala 47:23]
  reg [184:0] cache_data_751; // @[icache.scala 47:23]
  reg [184:0] cache_data_752; // @[icache.scala 47:23]
  reg [184:0] cache_data_753; // @[icache.scala 47:23]
  reg [184:0] cache_data_754; // @[icache.scala 47:23]
  reg [184:0] cache_data_755; // @[icache.scala 47:23]
  reg [184:0] cache_data_756; // @[icache.scala 47:23]
  reg [184:0] cache_data_757; // @[icache.scala 47:23]
  reg [184:0] cache_data_758; // @[icache.scala 47:23]
  reg [184:0] cache_data_759; // @[icache.scala 47:23]
  reg [184:0] cache_data_760; // @[icache.scala 47:23]
  reg [184:0] cache_data_761; // @[icache.scala 47:23]
  reg [184:0] cache_data_762; // @[icache.scala 47:23]
  reg [184:0] cache_data_763; // @[icache.scala 47:23]
  reg [184:0] cache_data_764; // @[icache.scala 47:23]
  reg [184:0] cache_data_765; // @[icache.scala 47:23]
  reg [184:0] cache_data_766; // @[icache.scala 47:23]
  reg [184:0] cache_data_767; // @[icache.scala 47:23]
  reg [184:0] cache_data_768; // @[icache.scala 47:23]
  reg [184:0] cache_data_769; // @[icache.scala 47:23]
  reg [184:0] cache_data_770; // @[icache.scala 47:23]
  reg [184:0] cache_data_771; // @[icache.scala 47:23]
  reg [184:0] cache_data_772; // @[icache.scala 47:23]
  reg [184:0] cache_data_773; // @[icache.scala 47:23]
  reg [184:0] cache_data_774; // @[icache.scala 47:23]
  reg [184:0] cache_data_775; // @[icache.scala 47:23]
  reg [184:0] cache_data_776; // @[icache.scala 47:23]
  reg [184:0] cache_data_777; // @[icache.scala 47:23]
  reg [184:0] cache_data_778; // @[icache.scala 47:23]
  reg [184:0] cache_data_779; // @[icache.scala 47:23]
  reg [184:0] cache_data_780; // @[icache.scala 47:23]
  reg [184:0] cache_data_781; // @[icache.scala 47:23]
  reg [184:0] cache_data_782; // @[icache.scala 47:23]
  reg [184:0] cache_data_783; // @[icache.scala 47:23]
  reg [184:0] cache_data_784; // @[icache.scala 47:23]
  reg [184:0] cache_data_785; // @[icache.scala 47:23]
  reg [184:0] cache_data_786; // @[icache.scala 47:23]
  reg [184:0] cache_data_787; // @[icache.scala 47:23]
  reg [184:0] cache_data_788; // @[icache.scala 47:23]
  reg [184:0] cache_data_789; // @[icache.scala 47:23]
  reg [184:0] cache_data_790; // @[icache.scala 47:23]
  reg [184:0] cache_data_791; // @[icache.scala 47:23]
  reg [184:0] cache_data_792; // @[icache.scala 47:23]
  reg [184:0] cache_data_793; // @[icache.scala 47:23]
  reg [184:0] cache_data_794; // @[icache.scala 47:23]
  reg [184:0] cache_data_795; // @[icache.scala 47:23]
  reg [184:0] cache_data_796; // @[icache.scala 47:23]
  reg [184:0] cache_data_797; // @[icache.scala 47:23]
  reg [184:0] cache_data_798; // @[icache.scala 47:23]
  reg [184:0] cache_data_799; // @[icache.scala 47:23]
  reg [184:0] cache_data_800; // @[icache.scala 47:23]
  reg [184:0] cache_data_801; // @[icache.scala 47:23]
  reg [184:0] cache_data_802; // @[icache.scala 47:23]
  reg [184:0] cache_data_803; // @[icache.scala 47:23]
  reg [184:0] cache_data_804; // @[icache.scala 47:23]
  reg [184:0] cache_data_805; // @[icache.scala 47:23]
  reg [184:0] cache_data_806; // @[icache.scala 47:23]
  reg [184:0] cache_data_807; // @[icache.scala 47:23]
  reg [184:0] cache_data_808; // @[icache.scala 47:23]
  reg [184:0] cache_data_809; // @[icache.scala 47:23]
  reg [184:0] cache_data_810; // @[icache.scala 47:23]
  reg [184:0] cache_data_811; // @[icache.scala 47:23]
  reg [184:0] cache_data_812; // @[icache.scala 47:23]
  reg [184:0] cache_data_813; // @[icache.scala 47:23]
  reg [184:0] cache_data_814; // @[icache.scala 47:23]
  reg [184:0] cache_data_815; // @[icache.scala 47:23]
  reg [184:0] cache_data_816; // @[icache.scala 47:23]
  reg [184:0] cache_data_817; // @[icache.scala 47:23]
  reg [184:0] cache_data_818; // @[icache.scala 47:23]
  reg [184:0] cache_data_819; // @[icache.scala 47:23]
  reg [184:0] cache_data_820; // @[icache.scala 47:23]
  reg [184:0] cache_data_821; // @[icache.scala 47:23]
  reg [184:0] cache_data_822; // @[icache.scala 47:23]
  reg [184:0] cache_data_823; // @[icache.scala 47:23]
  reg [184:0] cache_data_824; // @[icache.scala 47:23]
  reg [184:0] cache_data_825; // @[icache.scala 47:23]
  reg [184:0] cache_data_826; // @[icache.scala 47:23]
  reg [184:0] cache_data_827; // @[icache.scala 47:23]
  reg [184:0] cache_data_828; // @[icache.scala 47:23]
  reg [184:0] cache_data_829; // @[icache.scala 47:23]
  reg [184:0] cache_data_830; // @[icache.scala 47:23]
  reg [184:0] cache_data_831; // @[icache.scala 47:23]
  reg [184:0] cache_data_832; // @[icache.scala 47:23]
  reg [184:0] cache_data_833; // @[icache.scala 47:23]
  reg [184:0] cache_data_834; // @[icache.scala 47:23]
  reg [184:0] cache_data_835; // @[icache.scala 47:23]
  reg [184:0] cache_data_836; // @[icache.scala 47:23]
  reg [184:0] cache_data_837; // @[icache.scala 47:23]
  reg [184:0] cache_data_838; // @[icache.scala 47:23]
  reg [184:0] cache_data_839; // @[icache.scala 47:23]
  reg [184:0] cache_data_840; // @[icache.scala 47:23]
  reg [184:0] cache_data_841; // @[icache.scala 47:23]
  reg [184:0] cache_data_842; // @[icache.scala 47:23]
  reg [184:0] cache_data_843; // @[icache.scala 47:23]
  reg [184:0] cache_data_844; // @[icache.scala 47:23]
  reg [184:0] cache_data_845; // @[icache.scala 47:23]
  reg [184:0] cache_data_846; // @[icache.scala 47:23]
  reg [184:0] cache_data_847; // @[icache.scala 47:23]
  reg [184:0] cache_data_848; // @[icache.scala 47:23]
  reg [184:0] cache_data_849; // @[icache.scala 47:23]
  reg [184:0] cache_data_850; // @[icache.scala 47:23]
  reg [184:0] cache_data_851; // @[icache.scala 47:23]
  reg [184:0] cache_data_852; // @[icache.scala 47:23]
  reg [184:0] cache_data_853; // @[icache.scala 47:23]
  reg [184:0] cache_data_854; // @[icache.scala 47:23]
  reg [184:0] cache_data_855; // @[icache.scala 47:23]
  reg [184:0] cache_data_856; // @[icache.scala 47:23]
  reg [184:0] cache_data_857; // @[icache.scala 47:23]
  reg [184:0] cache_data_858; // @[icache.scala 47:23]
  reg [184:0] cache_data_859; // @[icache.scala 47:23]
  reg [184:0] cache_data_860; // @[icache.scala 47:23]
  reg [184:0] cache_data_861; // @[icache.scala 47:23]
  reg [184:0] cache_data_862; // @[icache.scala 47:23]
  reg [184:0] cache_data_863; // @[icache.scala 47:23]
  reg [184:0] cache_data_864; // @[icache.scala 47:23]
  reg [184:0] cache_data_865; // @[icache.scala 47:23]
  reg [184:0] cache_data_866; // @[icache.scala 47:23]
  reg [184:0] cache_data_867; // @[icache.scala 47:23]
  reg [184:0] cache_data_868; // @[icache.scala 47:23]
  reg [184:0] cache_data_869; // @[icache.scala 47:23]
  reg [184:0] cache_data_870; // @[icache.scala 47:23]
  reg [184:0] cache_data_871; // @[icache.scala 47:23]
  reg [184:0] cache_data_872; // @[icache.scala 47:23]
  reg [184:0] cache_data_873; // @[icache.scala 47:23]
  reg [184:0] cache_data_874; // @[icache.scala 47:23]
  reg [184:0] cache_data_875; // @[icache.scala 47:23]
  reg [184:0] cache_data_876; // @[icache.scala 47:23]
  reg [184:0] cache_data_877; // @[icache.scala 47:23]
  reg [184:0] cache_data_878; // @[icache.scala 47:23]
  reg [184:0] cache_data_879; // @[icache.scala 47:23]
  reg [184:0] cache_data_880; // @[icache.scala 47:23]
  reg [184:0] cache_data_881; // @[icache.scala 47:23]
  reg [184:0] cache_data_882; // @[icache.scala 47:23]
  reg [184:0] cache_data_883; // @[icache.scala 47:23]
  reg [184:0] cache_data_884; // @[icache.scala 47:23]
  reg [184:0] cache_data_885; // @[icache.scala 47:23]
  reg [184:0] cache_data_886; // @[icache.scala 47:23]
  reg [184:0] cache_data_887; // @[icache.scala 47:23]
  reg [184:0] cache_data_888; // @[icache.scala 47:23]
  reg [184:0] cache_data_889; // @[icache.scala 47:23]
  reg [184:0] cache_data_890; // @[icache.scala 47:23]
  reg [184:0] cache_data_891; // @[icache.scala 47:23]
  reg [184:0] cache_data_892; // @[icache.scala 47:23]
  reg [184:0] cache_data_893; // @[icache.scala 47:23]
  reg [184:0] cache_data_894; // @[icache.scala 47:23]
  reg [184:0] cache_data_895; // @[icache.scala 47:23]
  reg [184:0] cache_data_896; // @[icache.scala 47:23]
  reg [184:0] cache_data_897; // @[icache.scala 47:23]
  reg [184:0] cache_data_898; // @[icache.scala 47:23]
  reg [184:0] cache_data_899; // @[icache.scala 47:23]
  reg [184:0] cache_data_900; // @[icache.scala 47:23]
  reg [184:0] cache_data_901; // @[icache.scala 47:23]
  reg [184:0] cache_data_902; // @[icache.scala 47:23]
  reg [184:0] cache_data_903; // @[icache.scala 47:23]
  reg [184:0] cache_data_904; // @[icache.scala 47:23]
  reg [184:0] cache_data_905; // @[icache.scala 47:23]
  reg [184:0] cache_data_906; // @[icache.scala 47:23]
  reg [184:0] cache_data_907; // @[icache.scala 47:23]
  reg [184:0] cache_data_908; // @[icache.scala 47:23]
  reg [184:0] cache_data_909; // @[icache.scala 47:23]
  reg [184:0] cache_data_910; // @[icache.scala 47:23]
  reg [184:0] cache_data_911; // @[icache.scala 47:23]
  reg [184:0] cache_data_912; // @[icache.scala 47:23]
  reg [184:0] cache_data_913; // @[icache.scala 47:23]
  reg [184:0] cache_data_914; // @[icache.scala 47:23]
  reg [184:0] cache_data_915; // @[icache.scala 47:23]
  reg [184:0] cache_data_916; // @[icache.scala 47:23]
  reg [184:0] cache_data_917; // @[icache.scala 47:23]
  reg [184:0] cache_data_918; // @[icache.scala 47:23]
  reg [184:0] cache_data_919; // @[icache.scala 47:23]
  reg [184:0] cache_data_920; // @[icache.scala 47:23]
  reg [184:0] cache_data_921; // @[icache.scala 47:23]
  reg [184:0] cache_data_922; // @[icache.scala 47:23]
  reg [184:0] cache_data_923; // @[icache.scala 47:23]
  reg [184:0] cache_data_924; // @[icache.scala 47:23]
  reg [184:0] cache_data_925; // @[icache.scala 47:23]
  reg [184:0] cache_data_926; // @[icache.scala 47:23]
  reg [184:0] cache_data_927; // @[icache.scala 47:23]
  reg [184:0] cache_data_928; // @[icache.scala 47:23]
  reg [184:0] cache_data_929; // @[icache.scala 47:23]
  reg [184:0] cache_data_930; // @[icache.scala 47:23]
  reg [184:0] cache_data_931; // @[icache.scala 47:23]
  reg [184:0] cache_data_932; // @[icache.scala 47:23]
  reg [184:0] cache_data_933; // @[icache.scala 47:23]
  reg [184:0] cache_data_934; // @[icache.scala 47:23]
  reg [184:0] cache_data_935; // @[icache.scala 47:23]
  reg [184:0] cache_data_936; // @[icache.scala 47:23]
  reg [184:0] cache_data_937; // @[icache.scala 47:23]
  reg [184:0] cache_data_938; // @[icache.scala 47:23]
  reg [184:0] cache_data_939; // @[icache.scala 47:23]
  reg [184:0] cache_data_940; // @[icache.scala 47:23]
  reg [184:0] cache_data_941; // @[icache.scala 47:23]
  reg [184:0] cache_data_942; // @[icache.scala 47:23]
  reg [184:0] cache_data_943; // @[icache.scala 47:23]
  reg [184:0] cache_data_944; // @[icache.scala 47:23]
  reg [184:0] cache_data_945; // @[icache.scala 47:23]
  reg [184:0] cache_data_946; // @[icache.scala 47:23]
  reg [184:0] cache_data_947; // @[icache.scala 47:23]
  reg [184:0] cache_data_948; // @[icache.scala 47:23]
  reg [184:0] cache_data_949; // @[icache.scala 47:23]
  reg [184:0] cache_data_950; // @[icache.scala 47:23]
  reg [184:0] cache_data_951; // @[icache.scala 47:23]
  reg [184:0] cache_data_952; // @[icache.scala 47:23]
  reg [184:0] cache_data_953; // @[icache.scala 47:23]
  reg [184:0] cache_data_954; // @[icache.scala 47:23]
  reg [184:0] cache_data_955; // @[icache.scala 47:23]
  reg [184:0] cache_data_956; // @[icache.scala 47:23]
  reg [184:0] cache_data_957; // @[icache.scala 47:23]
  reg [184:0] cache_data_958; // @[icache.scala 47:23]
  reg [184:0] cache_data_959; // @[icache.scala 47:23]
  reg [184:0] cache_data_960; // @[icache.scala 47:23]
  reg [184:0] cache_data_961; // @[icache.scala 47:23]
  reg [184:0] cache_data_962; // @[icache.scala 47:23]
  reg [184:0] cache_data_963; // @[icache.scala 47:23]
  reg [184:0] cache_data_964; // @[icache.scala 47:23]
  reg [184:0] cache_data_965; // @[icache.scala 47:23]
  reg [184:0] cache_data_966; // @[icache.scala 47:23]
  reg [184:0] cache_data_967; // @[icache.scala 47:23]
  reg [184:0] cache_data_968; // @[icache.scala 47:23]
  reg [184:0] cache_data_969; // @[icache.scala 47:23]
  reg [184:0] cache_data_970; // @[icache.scala 47:23]
  reg [184:0] cache_data_971; // @[icache.scala 47:23]
  reg [184:0] cache_data_972; // @[icache.scala 47:23]
  reg [184:0] cache_data_973; // @[icache.scala 47:23]
  reg [184:0] cache_data_974; // @[icache.scala 47:23]
  reg [184:0] cache_data_975; // @[icache.scala 47:23]
  reg [184:0] cache_data_976; // @[icache.scala 47:23]
  reg [184:0] cache_data_977; // @[icache.scala 47:23]
  reg [184:0] cache_data_978; // @[icache.scala 47:23]
  reg [184:0] cache_data_979; // @[icache.scala 47:23]
  reg [184:0] cache_data_980; // @[icache.scala 47:23]
  reg [184:0] cache_data_981; // @[icache.scala 47:23]
  reg [184:0] cache_data_982; // @[icache.scala 47:23]
  reg [184:0] cache_data_983; // @[icache.scala 47:23]
  reg [184:0] cache_data_984; // @[icache.scala 47:23]
  reg [184:0] cache_data_985; // @[icache.scala 47:23]
  reg [184:0] cache_data_986; // @[icache.scala 47:23]
  reg [184:0] cache_data_987; // @[icache.scala 47:23]
  reg [184:0] cache_data_988; // @[icache.scala 47:23]
  reg [184:0] cache_data_989; // @[icache.scala 47:23]
  reg [184:0] cache_data_990; // @[icache.scala 47:23]
  reg [184:0] cache_data_991; // @[icache.scala 47:23]
  reg [184:0] cache_data_992; // @[icache.scala 47:23]
  reg [184:0] cache_data_993; // @[icache.scala 47:23]
  reg [184:0] cache_data_994; // @[icache.scala 47:23]
  reg [184:0] cache_data_995; // @[icache.scala 47:23]
  reg [184:0] cache_data_996; // @[icache.scala 47:23]
  reg [184:0] cache_data_997; // @[icache.scala 47:23]
  reg [184:0] cache_data_998; // @[icache.scala 47:23]
  reg [184:0] cache_data_999; // @[icache.scala 47:23]
  reg [184:0] cache_data_1000; // @[icache.scala 47:23]
  reg [184:0] cache_data_1001; // @[icache.scala 47:23]
  reg [184:0] cache_data_1002; // @[icache.scala 47:23]
  reg [184:0] cache_data_1003; // @[icache.scala 47:23]
  reg [184:0] cache_data_1004; // @[icache.scala 47:23]
  reg [184:0] cache_data_1005; // @[icache.scala 47:23]
  reg [184:0] cache_data_1006; // @[icache.scala 47:23]
  reg [184:0] cache_data_1007; // @[icache.scala 47:23]
  reg [184:0] cache_data_1008; // @[icache.scala 47:23]
  reg [184:0] cache_data_1009; // @[icache.scala 47:23]
  reg [184:0] cache_data_1010; // @[icache.scala 47:23]
  reg [184:0] cache_data_1011; // @[icache.scala 47:23]
  reg [184:0] cache_data_1012; // @[icache.scala 47:23]
  reg [184:0] cache_data_1013; // @[icache.scala 47:23]
  reg [184:0] cache_data_1014; // @[icache.scala 47:23]
  reg [184:0] cache_data_1015; // @[icache.scala 47:23]
  reg [184:0] cache_data_1016; // @[icache.scala 47:23]
  reg [184:0] cache_data_1017; // @[icache.scala 47:23]
  reg [184:0] cache_data_1018; // @[icache.scala 47:23]
  reg [184:0] cache_data_1019; // @[icache.scala 47:23]
  reg [184:0] cache_data_1020; // @[icache.scala 47:23]
  reg [184:0] cache_data_1021; // @[icache.scala 47:23]
  reg [184:0] cache_data_1022; // @[icache.scala 47:23]
  reg [184:0] cache_data_1023; // @[icache.scala 47:23]
  wire [184:0] _GEN_1 = 10'h1 == cpu_index ? cache_data_1 : cache_data_0; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_2 = 10'h2 == cpu_index ? cache_data_2 : _GEN_1; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_3 = 10'h3 == cpu_index ? cache_data_3 : _GEN_2; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_4 = 10'h4 == cpu_index ? cache_data_4 : _GEN_3; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_5 = 10'h5 == cpu_index ? cache_data_5 : _GEN_4; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_6 = 10'h6 == cpu_index ? cache_data_6 : _GEN_5; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_7 = 10'h7 == cpu_index ? cache_data_7 : _GEN_6; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_8 = 10'h8 == cpu_index ? cache_data_8 : _GEN_7; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_9 = 10'h9 == cpu_index ? cache_data_9 : _GEN_8; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_10 = 10'ha == cpu_index ? cache_data_10 : _GEN_9; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_11 = 10'hb == cpu_index ? cache_data_11 : _GEN_10; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_12 = 10'hc == cpu_index ? cache_data_12 : _GEN_11; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_13 = 10'hd == cpu_index ? cache_data_13 : _GEN_12; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_14 = 10'he == cpu_index ? cache_data_14 : _GEN_13; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_15 = 10'hf == cpu_index ? cache_data_15 : _GEN_14; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_16 = 10'h10 == cpu_index ? cache_data_16 : _GEN_15; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_17 = 10'h11 == cpu_index ? cache_data_17 : _GEN_16; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_18 = 10'h12 == cpu_index ? cache_data_18 : _GEN_17; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_19 = 10'h13 == cpu_index ? cache_data_19 : _GEN_18; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_20 = 10'h14 == cpu_index ? cache_data_20 : _GEN_19; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_21 = 10'h15 == cpu_index ? cache_data_21 : _GEN_20; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_22 = 10'h16 == cpu_index ? cache_data_22 : _GEN_21; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_23 = 10'h17 == cpu_index ? cache_data_23 : _GEN_22; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_24 = 10'h18 == cpu_index ? cache_data_24 : _GEN_23; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_25 = 10'h19 == cpu_index ? cache_data_25 : _GEN_24; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_26 = 10'h1a == cpu_index ? cache_data_26 : _GEN_25; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_27 = 10'h1b == cpu_index ? cache_data_27 : _GEN_26; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_28 = 10'h1c == cpu_index ? cache_data_28 : _GEN_27; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_29 = 10'h1d == cpu_index ? cache_data_29 : _GEN_28; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_30 = 10'h1e == cpu_index ? cache_data_30 : _GEN_29; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_31 = 10'h1f == cpu_index ? cache_data_31 : _GEN_30; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_32 = 10'h20 == cpu_index ? cache_data_32 : _GEN_31; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_33 = 10'h21 == cpu_index ? cache_data_33 : _GEN_32; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_34 = 10'h22 == cpu_index ? cache_data_34 : _GEN_33; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_35 = 10'h23 == cpu_index ? cache_data_35 : _GEN_34; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_36 = 10'h24 == cpu_index ? cache_data_36 : _GEN_35; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_37 = 10'h25 == cpu_index ? cache_data_37 : _GEN_36; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_38 = 10'h26 == cpu_index ? cache_data_38 : _GEN_37; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_39 = 10'h27 == cpu_index ? cache_data_39 : _GEN_38; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_40 = 10'h28 == cpu_index ? cache_data_40 : _GEN_39; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_41 = 10'h29 == cpu_index ? cache_data_41 : _GEN_40; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_42 = 10'h2a == cpu_index ? cache_data_42 : _GEN_41; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_43 = 10'h2b == cpu_index ? cache_data_43 : _GEN_42; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_44 = 10'h2c == cpu_index ? cache_data_44 : _GEN_43; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_45 = 10'h2d == cpu_index ? cache_data_45 : _GEN_44; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_46 = 10'h2e == cpu_index ? cache_data_46 : _GEN_45; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_47 = 10'h2f == cpu_index ? cache_data_47 : _GEN_46; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_48 = 10'h30 == cpu_index ? cache_data_48 : _GEN_47; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_49 = 10'h31 == cpu_index ? cache_data_49 : _GEN_48; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_50 = 10'h32 == cpu_index ? cache_data_50 : _GEN_49; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_51 = 10'h33 == cpu_index ? cache_data_51 : _GEN_50; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_52 = 10'h34 == cpu_index ? cache_data_52 : _GEN_51; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_53 = 10'h35 == cpu_index ? cache_data_53 : _GEN_52; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_54 = 10'h36 == cpu_index ? cache_data_54 : _GEN_53; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_55 = 10'h37 == cpu_index ? cache_data_55 : _GEN_54; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_56 = 10'h38 == cpu_index ? cache_data_56 : _GEN_55; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_57 = 10'h39 == cpu_index ? cache_data_57 : _GEN_56; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_58 = 10'h3a == cpu_index ? cache_data_58 : _GEN_57; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_59 = 10'h3b == cpu_index ? cache_data_59 : _GEN_58; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_60 = 10'h3c == cpu_index ? cache_data_60 : _GEN_59; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_61 = 10'h3d == cpu_index ? cache_data_61 : _GEN_60; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_62 = 10'h3e == cpu_index ? cache_data_62 : _GEN_61; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_63 = 10'h3f == cpu_index ? cache_data_63 : _GEN_62; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_64 = 10'h40 == cpu_index ? cache_data_64 : _GEN_63; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_65 = 10'h41 == cpu_index ? cache_data_65 : _GEN_64; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_66 = 10'h42 == cpu_index ? cache_data_66 : _GEN_65; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_67 = 10'h43 == cpu_index ? cache_data_67 : _GEN_66; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_68 = 10'h44 == cpu_index ? cache_data_68 : _GEN_67; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_69 = 10'h45 == cpu_index ? cache_data_69 : _GEN_68; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_70 = 10'h46 == cpu_index ? cache_data_70 : _GEN_69; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_71 = 10'h47 == cpu_index ? cache_data_71 : _GEN_70; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_72 = 10'h48 == cpu_index ? cache_data_72 : _GEN_71; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_73 = 10'h49 == cpu_index ? cache_data_73 : _GEN_72; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_74 = 10'h4a == cpu_index ? cache_data_74 : _GEN_73; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_75 = 10'h4b == cpu_index ? cache_data_75 : _GEN_74; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_76 = 10'h4c == cpu_index ? cache_data_76 : _GEN_75; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_77 = 10'h4d == cpu_index ? cache_data_77 : _GEN_76; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_78 = 10'h4e == cpu_index ? cache_data_78 : _GEN_77; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_79 = 10'h4f == cpu_index ? cache_data_79 : _GEN_78; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_80 = 10'h50 == cpu_index ? cache_data_80 : _GEN_79; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_81 = 10'h51 == cpu_index ? cache_data_81 : _GEN_80; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_82 = 10'h52 == cpu_index ? cache_data_82 : _GEN_81; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_83 = 10'h53 == cpu_index ? cache_data_83 : _GEN_82; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_84 = 10'h54 == cpu_index ? cache_data_84 : _GEN_83; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_85 = 10'h55 == cpu_index ? cache_data_85 : _GEN_84; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_86 = 10'h56 == cpu_index ? cache_data_86 : _GEN_85; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_87 = 10'h57 == cpu_index ? cache_data_87 : _GEN_86; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_88 = 10'h58 == cpu_index ? cache_data_88 : _GEN_87; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_89 = 10'h59 == cpu_index ? cache_data_89 : _GEN_88; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_90 = 10'h5a == cpu_index ? cache_data_90 : _GEN_89; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_91 = 10'h5b == cpu_index ? cache_data_91 : _GEN_90; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_92 = 10'h5c == cpu_index ? cache_data_92 : _GEN_91; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_93 = 10'h5d == cpu_index ? cache_data_93 : _GEN_92; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_94 = 10'h5e == cpu_index ? cache_data_94 : _GEN_93; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_95 = 10'h5f == cpu_index ? cache_data_95 : _GEN_94; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_96 = 10'h60 == cpu_index ? cache_data_96 : _GEN_95; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_97 = 10'h61 == cpu_index ? cache_data_97 : _GEN_96; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_98 = 10'h62 == cpu_index ? cache_data_98 : _GEN_97; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_99 = 10'h63 == cpu_index ? cache_data_99 : _GEN_98; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_100 = 10'h64 == cpu_index ? cache_data_100 : _GEN_99; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_101 = 10'h65 == cpu_index ? cache_data_101 : _GEN_100; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_102 = 10'h66 == cpu_index ? cache_data_102 : _GEN_101; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_103 = 10'h67 == cpu_index ? cache_data_103 : _GEN_102; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_104 = 10'h68 == cpu_index ? cache_data_104 : _GEN_103; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_105 = 10'h69 == cpu_index ? cache_data_105 : _GEN_104; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_106 = 10'h6a == cpu_index ? cache_data_106 : _GEN_105; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_107 = 10'h6b == cpu_index ? cache_data_107 : _GEN_106; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_108 = 10'h6c == cpu_index ? cache_data_108 : _GEN_107; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_109 = 10'h6d == cpu_index ? cache_data_109 : _GEN_108; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_110 = 10'h6e == cpu_index ? cache_data_110 : _GEN_109; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_111 = 10'h6f == cpu_index ? cache_data_111 : _GEN_110; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_112 = 10'h70 == cpu_index ? cache_data_112 : _GEN_111; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_113 = 10'h71 == cpu_index ? cache_data_113 : _GEN_112; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_114 = 10'h72 == cpu_index ? cache_data_114 : _GEN_113; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_115 = 10'h73 == cpu_index ? cache_data_115 : _GEN_114; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_116 = 10'h74 == cpu_index ? cache_data_116 : _GEN_115; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_117 = 10'h75 == cpu_index ? cache_data_117 : _GEN_116; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_118 = 10'h76 == cpu_index ? cache_data_118 : _GEN_117; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_119 = 10'h77 == cpu_index ? cache_data_119 : _GEN_118; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_120 = 10'h78 == cpu_index ? cache_data_120 : _GEN_119; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_121 = 10'h79 == cpu_index ? cache_data_121 : _GEN_120; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_122 = 10'h7a == cpu_index ? cache_data_122 : _GEN_121; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_123 = 10'h7b == cpu_index ? cache_data_123 : _GEN_122; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_124 = 10'h7c == cpu_index ? cache_data_124 : _GEN_123; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_125 = 10'h7d == cpu_index ? cache_data_125 : _GEN_124; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_126 = 10'h7e == cpu_index ? cache_data_126 : _GEN_125; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_127 = 10'h7f == cpu_index ? cache_data_127 : _GEN_126; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_128 = 10'h80 == cpu_index ? cache_data_128 : _GEN_127; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_129 = 10'h81 == cpu_index ? cache_data_129 : _GEN_128; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_130 = 10'h82 == cpu_index ? cache_data_130 : _GEN_129; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_131 = 10'h83 == cpu_index ? cache_data_131 : _GEN_130; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_132 = 10'h84 == cpu_index ? cache_data_132 : _GEN_131; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_133 = 10'h85 == cpu_index ? cache_data_133 : _GEN_132; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_134 = 10'h86 == cpu_index ? cache_data_134 : _GEN_133; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_135 = 10'h87 == cpu_index ? cache_data_135 : _GEN_134; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_136 = 10'h88 == cpu_index ? cache_data_136 : _GEN_135; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_137 = 10'h89 == cpu_index ? cache_data_137 : _GEN_136; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_138 = 10'h8a == cpu_index ? cache_data_138 : _GEN_137; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_139 = 10'h8b == cpu_index ? cache_data_139 : _GEN_138; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_140 = 10'h8c == cpu_index ? cache_data_140 : _GEN_139; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_141 = 10'h8d == cpu_index ? cache_data_141 : _GEN_140; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_142 = 10'h8e == cpu_index ? cache_data_142 : _GEN_141; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_143 = 10'h8f == cpu_index ? cache_data_143 : _GEN_142; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_144 = 10'h90 == cpu_index ? cache_data_144 : _GEN_143; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_145 = 10'h91 == cpu_index ? cache_data_145 : _GEN_144; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_146 = 10'h92 == cpu_index ? cache_data_146 : _GEN_145; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_147 = 10'h93 == cpu_index ? cache_data_147 : _GEN_146; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_148 = 10'h94 == cpu_index ? cache_data_148 : _GEN_147; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_149 = 10'h95 == cpu_index ? cache_data_149 : _GEN_148; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_150 = 10'h96 == cpu_index ? cache_data_150 : _GEN_149; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_151 = 10'h97 == cpu_index ? cache_data_151 : _GEN_150; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_152 = 10'h98 == cpu_index ? cache_data_152 : _GEN_151; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_153 = 10'h99 == cpu_index ? cache_data_153 : _GEN_152; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_154 = 10'h9a == cpu_index ? cache_data_154 : _GEN_153; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_155 = 10'h9b == cpu_index ? cache_data_155 : _GEN_154; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_156 = 10'h9c == cpu_index ? cache_data_156 : _GEN_155; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_157 = 10'h9d == cpu_index ? cache_data_157 : _GEN_156; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_158 = 10'h9e == cpu_index ? cache_data_158 : _GEN_157; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_159 = 10'h9f == cpu_index ? cache_data_159 : _GEN_158; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_160 = 10'ha0 == cpu_index ? cache_data_160 : _GEN_159; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_161 = 10'ha1 == cpu_index ? cache_data_161 : _GEN_160; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_162 = 10'ha2 == cpu_index ? cache_data_162 : _GEN_161; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_163 = 10'ha3 == cpu_index ? cache_data_163 : _GEN_162; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_164 = 10'ha4 == cpu_index ? cache_data_164 : _GEN_163; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_165 = 10'ha5 == cpu_index ? cache_data_165 : _GEN_164; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_166 = 10'ha6 == cpu_index ? cache_data_166 : _GEN_165; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_167 = 10'ha7 == cpu_index ? cache_data_167 : _GEN_166; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_168 = 10'ha8 == cpu_index ? cache_data_168 : _GEN_167; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_169 = 10'ha9 == cpu_index ? cache_data_169 : _GEN_168; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_170 = 10'haa == cpu_index ? cache_data_170 : _GEN_169; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_171 = 10'hab == cpu_index ? cache_data_171 : _GEN_170; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_172 = 10'hac == cpu_index ? cache_data_172 : _GEN_171; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_173 = 10'had == cpu_index ? cache_data_173 : _GEN_172; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_174 = 10'hae == cpu_index ? cache_data_174 : _GEN_173; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_175 = 10'haf == cpu_index ? cache_data_175 : _GEN_174; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_176 = 10'hb0 == cpu_index ? cache_data_176 : _GEN_175; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_177 = 10'hb1 == cpu_index ? cache_data_177 : _GEN_176; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_178 = 10'hb2 == cpu_index ? cache_data_178 : _GEN_177; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_179 = 10'hb3 == cpu_index ? cache_data_179 : _GEN_178; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_180 = 10'hb4 == cpu_index ? cache_data_180 : _GEN_179; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_181 = 10'hb5 == cpu_index ? cache_data_181 : _GEN_180; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_182 = 10'hb6 == cpu_index ? cache_data_182 : _GEN_181; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_183 = 10'hb7 == cpu_index ? cache_data_183 : _GEN_182; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_184 = 10'hb8 == cpu_index ? cache_data_184 : _GEN_183; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_185 = 10'hb9 == cpu_index ? cache_data_185 : _GEN_184; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_186 = 10'hba == cpu_index ? cache_data_186 : _GEN_185; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_187 = 10'hbb == cpu_index ? cache_data_187 : _GEN_186; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_188 = 10'hbc == cpu_index ? cache_data_188 : _GEN_187; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_189 = 10'hbd == cpu_index ? cache_data_189 : _GEN_188; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_190 = 10'hbe == cpu_index ? cache_data_190 : _GEN_189; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_191 = 10'hbf == cpu_index ? cache_data_191 : _GEN_190; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_192 = 10'hc0 == cpu_index ? cache_data_192 : _GEN_191; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_193 = 10'hc1 == cpu_index ? cache_data_193 : _GEN_192; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_194 = 10'hc2 == cpu_index ? cache_data_194 : _GEN_193; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_195 = 10'hc3 == cpu_index ? cache_data_195 : _GEN_194; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_196 = 10'hc4 == cpu_index ? cache_data_196 : _GEN_195; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_197 = 10'hc5 == cpu_index ? cache_data_197 : _GEN_196; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_198 = 10'hc6 == cpu_index ? cache_data_198 : _GEN_197; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_199 = 10'hc7 == cpu_index ? cache_data_199 : _GEN_198; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_200 = 10'hc8 == cpu_index ? cache_data_200 : _GEN_199; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_201 = 10'hc9 == cpu_index ? cache_data_201 : _GEN_200; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_202 = 10'hca == cpu_index ? cache_data_202 : _GEN_201; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_203 = 10'hcb == cpu_index ? cache_data_203 : _GEN_202; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_204 = 10'hcc == cpu_index ? cache_data_204 : _GEN_203; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_205 = 10'hcd == cpu_index ? cache_data_205 : _GEN_204; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_206 = 10'hce == cpu_index ? cache_data_206 : _GEN_205; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_207 = 10'hcf == cpu_index ? cache_data_207 : _GEN_206; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_208 = 10'hd0 == cpu_index ? cache_data_208 : _GEN_207; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_209 = 10'hd1 == cpu_index ? cache_data_209 : _GEN_208; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_210 = 10'hd2 == cpu_index ? cache_data_210 : _GEN_209; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_211 = 10'hd3 == cpu_index ? cache_data_211 : _GEN_210; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_212 = 10'hd4 == cpu_index ? cache_data_212 : _GEN_211; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_213 = 10'hd5 == cpu_index ? cache_data_213 : _GEN_212; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_214 = 10'hd6 == cpu_index ? cache_data_214 : _GEN_213; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_215 = 10'hd7 == cpu_index ? cache_data_215 : _GEN_214; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_216 = 10'hd8 == cpu_index ? cache_data_216 : _GEN_215; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_217 = 10'hd9 == cpu_index ? cache_data_217 : _GEN_216; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_218 = 10'hda == cpu_index ? cache_data_218 : _GEN_217; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_219 = 10'hdb == cpu_index ? cache_data_219 : _GEN_218; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_220 = 10'hdc == cpu_index ? cache_data_220 : _GEN_219; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_221 = 10'hdd == cpu_index ? cache_data_221 : _GEN_220; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_222 = 10'hde == cpu_index ? cache_data_222 : _GEN_221; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_223 = 10'hdf == cpu_index ? cache_data_223 : _GEN_222; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_224 = 10'he0 == cpu_index ? cache_data_224 : _GEN_223; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_225 = 10'he1 == cpu_index ? cache_data_225 : _GEN_224; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_226 = 10'he2 == cpu_index ? cache_data_226 : _GEN_225; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_227 = 10'he3 == cpu_index ? cache_data_227 : _GEN_226; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_228 = 10'he4 == cpu_index ? cache_data_228 : _GEN_227; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_229 = 10'he5 == cpu_index ? cache_data_229 : _GEN_228; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_230 = 10'he6 == cpu_index ? cache_data_230 : _GEN_229; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_231 = 10'he7 == cpu_index ? cache_data_231 : _GEN_230; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_232 = 10'he8 == cpu_index ? cache_data_232 : _GEN_231; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_233 = 10'he9 == cpu_index ? cache_data_233 : _GEN_232; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_234 = 10'hea == cpu_index ? cache_data_234 : _GEN_233; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_235 = 10'heb == cpu_index ? cache_data_235 : _GEN_234; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_236 = 10'hec == cpu_index ? cache_data_236 : _GEN_235; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_237 = 10'hed == cpu_index ? cache_data_237 : _GEN_236; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_238 = 10'hee == cpu_index ? cache_data_238 : _GEN_237; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_239 = 10'hef == cpu_index ? cache_data_239 : _GEN_238; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_240 = 10'hf0 == cpu_index ? cache_data_240 : _GEN_239; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_241 = 10'hf1 == cpu_index ? cache_data_241 : _GEN_240; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_242 = 10'hf2 == cpu_index ? cache_data_242 : _GEN_241; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_243 = 10'hf3 == cpu_index ? cache_data_243 : _GEN_242; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_244 = 10'hf4 == cpu_index ? cache_data_244 : _GEN_243; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_245 = 10'hf5 == cpu_index ? cache_data_245 : _GEN_244; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_246 = 10'hf6 == cpu_index ? cache_data_246 : _GEN_245; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_247 = 10'hf7 == cpu_index ? cache_data_247 : _GEN_246; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_248 = 10'hf8 == cpu_index ? cache_data_248 : _GEN_247; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_249 = 10'hf9 == cpu_index ? cache_data_249 : _GEN_248; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_250 = 10'hfa == cpu_index ? cache_data_250 : _GEN_249; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_251 = 10'hfb == cpu_index ? cache_data_251 : _GEN_250; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_252 = 10'hfc == cpu_index ? cache_data_252 : _GEN_251; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_253 = 10'hfd == cpu_index ? cache_data_253 : _GEN_252; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_254 = 10'hfe == cpu_index ? cache_data_254 : _GEN_253; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_255 = 10'hff == cpu_index ? cache_data_255 : _GEN_254; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_256 = 10'h100 == cpu_index ? cache_data_256 : _GEN_255; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_257 = 10'h101 == cpu_index ? cache_data_257 : _GEN_256; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_258 = 10'h102 == cpu_index ? cache_data_258 : _GEN_257; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_259 = 10'h103 == cpu_index ? cache_data_259 : _GEN_258; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_260 = 10'h104 == cpu_index ? cache_data_260 : _GEN_259; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_261 = 10'h105 == cpu_index ? cache_data_261 : _GEN_260; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_262 = 10'h106 == cpu_index ? cache_data_262 : _GEN_261; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_263 = 10'h107 == cpu_index ? cache_data_263 : _GEN_262; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_264 = 10'h108 == cpu_index ? cache_data_264 : _GEN_263; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_265 = 10'h109 == cpu_index ? cache_data_265 : _GEN_264; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_266 = 10'h10a == cpu_index ? cache_data_266 : _GEN_265; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_267 = 10'h10b == cpu_index ? cache_data_267 : _GEN_266; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_268 = 10'h10c == cpu_index ? cache_data_268 : _GEN_267; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_269 = 10'h10d == cpu_index ? cache_data_269 : _GEN_268; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_270 = 10'h10e == cpu_index ? cache_data_270 : _GEN_269; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_271 = 10'h10f == cpu_index ? cache_data_271 : _GEN_270; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_272 = 10'h110 == cpu_index ? cache_data_272 : _GEN_271; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_273 = 10'h111 == cpu_index ? cache_data_273 : _GEN_272; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_274 = 10'h112 == cpu_index ? cache_data_274 : _GEN_273; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_275 = 10'h113 == cpu_index ? cache_data_275 : _GEN_274; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_276 = 10'h114 == cpu_index ? cache_data_276 : _GEN_275; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_277 = 10'h115 == cpu_index ? cache_data_277 : _GEN_276; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_278 = 10'h116 == cpu_index ? cache_data_278 : _GEN_277; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_279 = 10'h117 == cpu_index ? cache_data_279 : _GEN_278; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_280 = 10'h118 == cpu_index ? cache_data_280 : _GEN_279; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_281 = 10'h119 == cpu_index ? cache_data_281 : _GEN_280; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_282 = 10'h11a == cpu_index ? cache_data_282 : _GEN_281; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_283 = 10'h11b == cpu_index ? cache_data_283 : _GEN_282; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_284 = 10'h11c == cpu_index ? cache_data_284 : _GEN_283; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_285 = 10'h11d == cpu_index ? cache_data_285 : _GEN_284; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_286 = 10'h11e == cpu_index ? cache_data_286 : _GEN_285; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_287 = 10'h11f == cpu_index ? cache_data_287 : _GEN_286; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_288 = 10'h120 == cpu_index ? cache_data_288 : _GEN_287; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_289 = 10'h121 == cpu_index ? cache_data_289 : _GEN_288; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_290 = 10'h122 == cpu_index ? cache_data_290 : _GEN_289; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_291 = 10'h123 == cpu_index ? cache_data_291 : _GEN_290; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_292 = 10'h124 == cpu_index ? cache_data_292 : _GEN_291; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_293 = 10'h125 == cpu_index ? cache_data_293 : _GEN_292; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_294 = 10'h126 == cpu_index ? cache_data_294 : _GEN_293; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_295 = 10'h127 == cpu_index ? cache_data_295 : _GEN_294; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_296 = 10'h128 == cpu_index ? cache_data_296 : _GEN_295; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_297 = 10'h129 == cpu_index ? cache_data_297 : _GEN_296; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_298 = 10'h12a == cpu_index ? cache_data_298 : _GEN_297; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_299 = 10'h12b == cpu_index ? cache_data_299 : _GEN_298; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_300 = 10'h12c == cpu_index ? cache_data_300 : _GEN_299; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_301 = 10'h12d == cpu_index ? cache_data_301 : _GEN_300; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_302 = 10'h12e == cpu_index ? cache_data_302 : _GEN_301; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_303 = 10'h12f == cpu_index ? cache_data_303 : _GEN_302; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_304 = 10'h130 == cpu_index ? cache_data_304 : _GEN_303; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_305 = 10'h131 == cpu_index ? cache_data_305 : _GEN_304; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_306 = 10'h132 == cpu_index ? cache_data_306 : _GEN_305; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_307 = 10'h133 == cpu_index ? cache_data_307 : _GEN_306; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_308 = 10'h134 == cpu_index ? cache_data_308 : _GEN_307; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_309 = 10'h135 == cpu_index ? cache_data_309 : _GEN_308; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_310 = 10'h136 == cpu_index ? cache_data_310 : _GEN_309; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_311 = 10'h137 == cpu_index ? cache_data_311 : _GEN_310; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_312 = 10'h138 == cpu_index ? cache_data_312 : _GEN_311; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_313 = 10'h139 == cpu_index ? cache_data_313 : _GEN_312; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_314 = 10'h13a == cpu_index ? cache_data_314 : _GEN_313; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_315 = 10'h13b == cpu_index ? cache_data_315 : _GEN_314; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_316 = 10'h13c == cpu_index ? cache_data_316 : _GEN_315; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_317 = 10'h13d == cpu_index ? cache_data_317 : _GEN_316; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_318 = 10'h13e == cpu_index ? cache_data_318 : _GEN_317; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_319 = 10'h13f == cpu_index ? cache_data_319 : _GEN_318; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_320 = 10'h140 == cpu_index ? cache_data_320 : _GEN_319; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_321 = 10'h141 == cpu_index ? cache_data_321 : _GEN_320; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_322 = 10'h142 == cpu_index ? cache_data_322 : _GEN_321; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_323 = 10'h143 == cpu_index ? cache_data_323 : _GEN_322; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_324 = 10'h144 == cpu_index ? cache_data_324 : _GEN_323; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_325 = 10'h145 == cpu_index ? cache_data_325 : _GEN_324; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_326 = 10'h146 == cpu_index ? cache_data_326 : _GEN_325; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_327 = 10'h147 == cpu_index ? cache_data_327 : _GEN_326; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_328 = 10'h148 == cpu_index ? cache_data_328 : _GEN_327; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_329 = 10'h149 == cpu_index ? cache_data_329 : _GEN_328; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_330 = 10'h14a == cpu_index ? cache_data_330 : _GEN_329; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_331 = 10'h14b == cpu_index ? cache_data_331 : _GEN_330; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_332 = 10'h14c == cpu_index ? cache_data_332 : _GEN_331; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_333 = 10'h14d == cpu_index ? cache_data_333 : _GEN_332; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_334 = 10'h14e == cpu_index ? cache_data_334 : _GEN_333; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_335 = 10'h14f == cpu_index ? cache_data_335 : _GEN_334; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_336 = 10'h150 == cpu_index ? cache_data_336 : _GEN_335; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_337 = 10'h151 == cpu_index ? cache_data_337 : _GEN_336; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_338 = 10'h152 == cpu_index ? cache_data_338 : _GEN_337; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_339 = 10'h153 == cpu_index ? cache_data_339 : _GEN_338; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_340 = 10'h154 == cpu_index ? cache_data_340 : _GEN_339; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_341 = 10'h155 == cpu_index ? cache_data_341 : _GEN_340; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_342 = 10'h156 == cpu_index ? cache_data_342 : _GEN_341; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_343 = 10'h157 == cpu_index ? cache_data_343 : _GEN_342; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_344 = 10'h158 == cpu_index ? cache_data_344 : _GEN_343; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_345 = 10'h159 == cpu_index ? cache_data_345 : _GEN_344; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_346 = 10'h15a == cpu_index ? cache_data_346 : _GEN_345; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_347 = 10'h15b == cpu_index ? cache_data_347 : _GEN_346; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_348 = 10'h15c == cpu_index ? cache_data_348 : _GEN_347; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_349 = 10'h15d == cpu_index ? cache_data_349 : _GEN_348; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_350 = 10'h15e == cpu_index ? cache_data_350 : _GEN_349; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_351 = 10'h15f == cpu_index ? cache_data_351 : _GEN_350; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_352 = 10'h160 == cpu_index ? cache_data_352 : _GEN_351; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_353 = 10'h161 == cpu_index ? cache_data_353 : _GEN_352; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_354 = 10'h162 == cpu_index ? cache_data_354 : _GEN_353; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_355 = 10'h163 == cpu_index ? cache_data_355 : _GEN_354; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_356 = 10'h164 == cpu_index ? cache_data_356 : _GEN_355; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_357 = 10'h165 == cpu_index ? cache_data_357 : _GEN_356; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_358 = 10'h166 == cpu_index ? cache_data_358 : _GEN_357; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_359 = 10'h167 == cpu_index ? cache_data_359 : _GEN_358; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_360 = 10'h168 == cpu_index ? cache_data_360 : _GEN_359; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_361 = 10'h169 == cpu_index ? cache_data_361 : _GEN_360; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_362 = 10'h16a == cpu_index ? cache_data_362 : _GEN_361; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_363 = 10'h16b == cpu_index ? cache_data_363 : _GEN_362; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_364 = 10'h16c == cpu_index ? cache_data_364 : _GEN_363; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_365 = 10'h16d == cpu_index ? cache_data_365 : _GEN_364; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_366 = 10'h16e == cpu_index ? cache_data_366 : _GEN_365; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_367 = 10'h16f == cpu_index ? cache_data_367 : _GEN_366; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_368 = 10'h170 == cpu_index ? cache_data_368 : _GEN_367; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_369 = 10'h171 == cpu_index ? cache_data_369 : _GEN_368; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_370 = 10'h172 == cpu_index ? cache_data_370 : _GEN_369; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_371 = 10'h173 == cpu_index ? cache_data_371 : _GEN_370; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_372 = 10'h174 == cpu_index ? cache_data_372 : _GEN_371; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_373 = 10'h175 == cpu_index ? cache_data_373 : _GEN_372; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_374 = 10'h176 == cpu_index ? cache_data_374 : _GEN_373; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_375 = 10'h177 == cpu_index ? cache_data_375 : _GEN_374; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_376 = 10'h178 == cpu_index ? cache_data_376 : _GEN_375; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_377 = 10'h179 == cpu_index ? cache_data_377 : _GEN_376; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_378 = 10'h17a == cpu_index ? cache_data_378 : _GEN_377; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_379 = 10'h17b == cpu_index ? cache_data_379 : _GEN_378; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_380 = 10'h17c == cpu_index ? cache_data_380 : _GEN_379; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_381 = 10'h17d == cpu_index ? cache_data_381 : _GEN_380; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_382 = 10'h17e == cpu_index ? cache_data_382 : _GEN_381; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_383 = 10'h17f == cpu_index ? cache_data_383 : _GEN_382; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_384 = 10'h180 == cpu_index ? cache_data_384 : _GEN_383; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_385 = 10'h181 == cpu_index ? cache_data_385 : _GEN_384; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_386 = 10'h182 == cpu_index ? cache_data_386 : _GEN_385; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_387 = 10'h183 == cpu_index ? cache_data_387 : _GEN_386; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_388 = 10'h184 == cpu_index ? cache_data_388 : _GEN_387; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_389 = 10'h185 == cpu_index ? cache_data_389 : _GEN_388; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_390 = 10'h186 == cpu_index ? cache_data_390 : _GEN_389; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_391 = 10'h187 == cpu_index ? cache_data_391 : _GEN_390; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_392 = 10'h188 == cpu_index ? cache_data_392 : _GEN_391; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_393 = 10'h189 == cpu_index ? cache_data_393 : _GEN_392; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_394 = 10'h18a == cpu_index ? cache_data_394 : _GEN_393; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_395 = 10'h18b == cpu_index ? cache_data_395 : _GEN_394; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_396 = 10'h18c == cpu_index ? cache_data_396 : _GEN_395; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_397 = 10'h18d == cpu_index ? cache_data_397 : _GEN_396; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_398 = 10'h18e == cpu_index ? cache_data_398 : _GEN_397; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_399 = 10'h18f == cpu_index ? cache_data_399 : _GEN_398; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_400 = 10'h190 == cpu_index ? cache_data_400 : _GEN_399; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_401 = 10'h191 == cpu_index ? cache_data_401 : _GEN_400; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_402 = 10'h192 == cpu_index ? cache_data_402 : _GEN_401; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_403 = 10'h193 == cpu_index ? cache_data_403 : _GEN_402; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_404 = 10'h194 == cpu_index ? cache_data_404 : _GEN_403; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_405 = 10'h195 == cpu_index ? cache_data_405 : _GEN_404; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_406 = 10'h196 == cpu_index ? cache_data_406 : _GEN_405; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_407 = 10'h197 == cpu_index ? cache_data_407 : _GEN_406; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_408 = 10'h198 == cpu_index ? cache_data_408 : _GEN_407; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_409 = 10'h199 == cpu_index ? cache_data_409 : _GEN_408; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_410 = 10'h19a == cpu_index ? cache_data_410 : _GEN_409; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_411 = 10'h19b == cpu_index ? cache_data_411 : _GEN_410; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_412 = 10'h19c == cpu_index ? cache_data_412 : _GEN_411; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_413 = 10'h19d == cpu_index ? cache_data_413 : _GEN_412; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_414 = 10'h19e == cpu_index ? cache_data_414 : _GEN_413; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_415 = 10'h19f == cpu_index ? cache_data_415 : _GEN_414; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_416 = 10'h1a0 == cpu_index ? cache_data_416 : _GEN_415; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_417 = 10'h1a1 == cpu_index ? cache_data_417 : _GEN_416; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_418 = 10'h1a2 == cpu_index ? cache_data_418 : _GEN_417; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_419 = 10'h1a3 == cpu_index ? cache_data_419 : _GEN_418; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_420 = 10'h1a4 == cpu_index ? cache_data_420 : _GEN_419; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_421 = 10'h1a5 == cpu_index ? cache_data_421 : _GEN_420; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_422 = 10'h1a6 == cpu_index ? cache_data_422 : _GEN_421; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_423 = 10'h1a7 == cpu_index ? cache_data_423 : _GEN_422; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_424 = 10'h1a8 == cpu_index ? cache_data_424 : _GEN_423; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_425 = 10'h1a9 == cpu_index ? cache_data_425 : _GEN_424; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_426 = 10'h1aa == cpu_index ? cache_data_426 : _GEN_425; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_427 = 10'h1ab == cpu_index ? cache_data_427 : _GEN_426; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_428 = 10'h1ac == cpu_index ? cache_data_428 : _GEN_427; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_429 = 10'h1ad == cpu_index ? cache_data_429 : _GEN_428; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_430 = 10'h1ae == cpu_index ? cache_data_430 : _GEN_429; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_431 = 10'h1af == cpu_index ? cache_data_431 : _GEN_430; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_432 = 10'h1b0 == cpu_index ? cache_data_432 : _GEN_431; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_433 = 10'h1b1 == cpu_index ? cache_data_433 : _GEN_432; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_434 = 10'h1b2 == cpu_index ? cache_data_434 : _GEN_433; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_435 = 10'h1b3 == cpu_index ? cache_data_435 : _GEN_434; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_436 = 10'h1b4 == cpu_index ? cache_data_436 : _GEN_435; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_437 = 10'h1b5 == cpu_index ? cache_data_437 : _GEN_436; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_438 = 10'h1b6 == cpu_index ? cache_data_438 : _GEN_437; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_439 = 10'h1b7 == cpu_index ? cache_data_439 : _GEN_438; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_440 = 10'h1b8 == cpu_index ? cache_data_440 : _GEN_439; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_441 = 10'h1b9 == cpu_index ? cache_data_441 : _GEN_440; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_442 = 10'h1ba == cpu_index ? cache_data_442 : _GEN_441; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_443 = 10'h1bb == cpu_index ? cache_data_443 : _GEN_442; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_444 = 10'h1bc == cpu_index ? cache_data_444 : _GEN_443; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_445 = 10'h1bd == cpu_index ? cache_data_445 : _GEN_444; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_446 = 10'h1be == cpu_index ? cache_data_446 : _GEN_445; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_447 = 10'h1bf == cpu_index ? cache_data_447 : _GEN_446; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_448 = 10'h1c0 == cpu_index ? cache_data_448 : _GEN_447; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_449 = 10'h1c1 == cpu_index ? cache_data_449 : _GEN_448; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_450 = 10'h1c2 == cpu_index ? cache_data_450 : _GEN_449; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_451 = 10'h1c3 == cpu_index ? cache_data_451 : _GEN_450; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_452 = 10'h1c4 == cpu_index ? cache_data_452 : _GEN_451; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_453 = 10'h1c5 == cpu_index ? cache_data_453 : _GEN_452; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_454 = 10'h1c6 == cpu_index ? cache_data_454 : _GEN_453; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_455 = 10'h1c7 == cpu_index ? cache_data_455 : _GEN_454; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_456 = 10'h1c8 == cpu_index ? cache_data_456 : _GEN_455; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_457 = 10'h1c9 == cpu_index ? cache_data_457 : _GEN_456; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_458 = 10'h1ca == cpu_index ? cache_data_458 : _GEN_457; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_459 = 10'h1cb == cpu_index ? cache_data_459 : _GEN_458; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_460 = 10'h1cc == cpu_index ? cache_data_460 : _GEN_459; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_461 = 10'h1cd == cpu_index ? cache_data_461 : _GEN_460; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_462 = 10'h1ce == cpu_index ? cache_data_462 : _GEN_461; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_463 = 10'h1cf == cpu_index ? cache_data_463 : _GEN_462; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_464 = 10'h1d0 == cpu_index ? cache_data_464 : _GEN_463; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_465 = 10'h1d1 == cpu_index ? cache_data_465 : _GEN_464; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_466 = 10'h1d2 == cpu_index ? cache_data_466 : _GEN_465; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_467 = 10'h1d3 == cpu_index ? cache_data_467 : _GEN_466; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_468 = 10'h1d4 == cpu_index ? cache_data_468 : _GEN_467; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_469 = 10'h1d5 == cpu_index ? cache_data_469 : _GEN_468; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_470 = 10'h1d6 == cpu_index ? cache_data_470 : _GEN_469; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_471 = 10'h1d7 == cpu_index ? cache_data_471 : _GEN_470; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_472 = 10'h1d8 == cpu_index ? cache_data_472 : _GEN_471; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_473 = 10'h1d9 == cpu_index ? cache_data_473 : _GEN_472; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_474 = 10'h1da == cpu_index ? cache_data_474 : _GEN_473; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_475 = 10'h1db == cpu_index ? cache_data_475 : _GEN_474; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_476 = 10'h1dc == cpu_index ? cache_data_476 : _GEN_475; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_477 = 10'h1dd == cpu_index ? cache_data_477 : _GEN_476; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_478 = 10'h1de == cpu_index ? cache_data_478 : _GEN_477; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_479 = 10'h1df == cpu_index ? cache_data_479 : _GEN_478; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_480 = 10'h1e0 == cpu_index ? cache_data_480 : _GEN_479; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_481 = 10'h1e1 == cpu_index ? cache_data_481 : _GEN_480; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_482 = 10'h1e2 == cpu_index ? cache_data_482 : _GEN_481; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_483 = 10'h1e3 == cpu_index ? cache_data_483 : _GEN_482; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_484 = 10'h1e4 == cpu_index ? cache_data_484 : _GEN_483; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_485 = 10'h1e5 == cpu_index ? cache_data_485 : _GEN_484; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_486 = 10'h1e6 == cpu_index ? cache_data_486 : _GEN_485; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_487 = 10'h1e7 == cpu_index ? cache_data_487 : _GEN_486; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_488 = 10'h1e8 == cpu_index ? cache_data_488 : _GEN_487; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_489 = 10'h1e9 == cpu_index ? cache_data_489 : _GEN_488; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_490 = 10'h1ea == cpu_index ? cache_data_490 : _GEN_489; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_491 = 10'h1eb == cpu_index ? cache_data_491 : _GEN_490; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_492 = 10'h1ec == cpu_index ? cache_data_492 : _GEN_491; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_493 = 10'h1ed == cpu_index ? cache_data_493 : _GEN_492; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_494 = 10'h1ee == cpu_index ? cache_data_494 : _GEN_493; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_495 = 10'h1ef == cpu_index ? cache_data_495 : _GEN_494; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_496 = 10'h1f0 == cpu_index ? cache_data_496 : _GEN_495; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_497 = 10'h1f1 == cpu_index ? cache_data_497 : _GEN_496; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_498 = 10'h1f2 == cpu_index ? cache_data_498 : _GEN_497; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_499 = 10'h1f3 == cpu_index ? cache_data_499 : _GEN_498; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_500 = 10'h1f4 == cpu_index ? cache_data_500 : _GEN_499; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_501 = 10'h1f5 == cpu_index ? cache_data_501 : _GEN_500; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_502 = 10'h1f6 == cpu_index ? cache_data_502 : _GEN_501; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_503 = 10'h1f7 == cpu_index ? cache_data_503 : _GEN_502; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_504 = 10'h1f8 == cpu_index ? cache_data_504 : _GEN_503; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_505 = 10'h1f9 == cpu_index ? cache_data_505 : _GEN_504; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_506 = 10'h1fa == cpu_index ? cache_data_506 : _GEN_505; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_507 = 10'h1fb == cpu_index ? cache_data_507 : _GEN_506; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_508 = 10'h1fc == cpu_index ? cache_data_508 : _GEN_507; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_509 = 10'h1fd == cpu_index ? cache_data_509 : _GEN_508; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_510 = 10'h1fe == cpu_index ? cache_data_510 : _GEN_509; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_511 = 10'h1ff == cpu_index ? cache_data_511 : _GEN_510; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_512 = 10'h200 == cpu_index ? cache_data_512 : _GEN_511; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_513 = 10'h201 == cpu_index ? cache_data_513 : _GEN_512; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_514 = 10'h202 == cpu_index ? cache_data_514 : _GEN_513; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_515 = 10'h203 == cpu_index ? cache_data_515 : _GEN_514; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_516 = 10'h204 == cpu_index ? cache_data_516 : _GEN_515; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_517 = 10'h205 == cpu_index ? cache_data_517 : _GEN_516; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_518 = 10'h206 == cpu_index ? cache_data_518 : _GEN_517; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_519 = 10'h207 == cpu_index ? cache_data_519 : _GEN_518; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_520 = 10'h208 == cpu_index ? cache_data_520 : _GEN_519; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_521 = 10'h209 == cpu_index ? cache_data_521 : _GEN_520; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_522 = 10'h20a == cpu_index ? cache_data_522 : _GEN_521; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_523 = 10'h20b == cpu_index ? cache_data_523 : _GEN_522; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_524 = 10'h20c == cpu_index ? cache_data_524 : _GEN_523; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_525 = 10'h20d == cpu_index ? cache_data_525 : _GEN_524; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_526 = 10'h20e == cpu_index ? cache_data_526 : _GEN_525; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_527 = 10'h20f == cpu_index ? cache_data_527 : _GEN_526; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_528 = 10'h210 == cpu_index ? cache_data_528 : _GEN_527; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_529 = 10'h211 == cpu_index ? cache_data_529 : _GEN_528; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_530 = 10'h212 == cpu_index ? cache_data_530 : _GEN_529; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_531 = 10'h213 == cpu_index ? cache_data_531 : _GEN_530; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_532 = 10'h214 == cpu_index ? cache_data_532 : _GEN_531; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_533 = 10'h215 == cpu_index ? cache_data_533 : _GEN_532; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_534 = 10'h216 == cpu_index ? cache_data_534 : _GEN_533; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_535 = 10'h217 == cpu_index ? cache_data_535 : _GEN_534; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_536 = 10'h218 == cpu_index ? cache_data_536 : _GEN_535; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_537 = 10'h219 == cpu_index ? cache_data_537 : _GEN_536; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_538 = 10'h21a == cpu_index ? cache_data_538 : _GEN_537; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_539 = 10'h21b == cpu_index ? cache_data_539 : _GEN_538; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_540 = 10'h21c == cpu_index ? cache_data_540 : _GEN_539; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_541 = 10'h21d == cpu_index ? cache_data_541 : _GEN_540; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_542 = 10'h21e == cpu_index ? cache_data_542 : _GEN_541; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_543 = 10'h21f == cpu_index ? cache_data_543 : _GEN_542; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_544 = 10'h220 == cpu_index ? cache_data_544 : _GEN_543; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_545 = 10'h221 == cpu_index ? cache_data_545 : _GEN_544; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_546 = 10'h222 == cpu_index ? cache_data_546 : _GEN_545; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_547 = 10'h223 == cpu_index ? cache_data_547 : _GEN_546; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_548 = 10'h224 == cpu_index ? cache_data_548 : _GEN_547; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_549 = 10'h225 == cpu_index ? cache_data_549 : _GEN_548; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_550 = 10'h226 == cpu_index ? cache_data_550 : _GEN_549; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_551 = 10'h227 == cpu_index ? cache_data_551 : _GEN_550; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_552 = 10'h228 == cpu_index ? cache_data_552 : _GEN_551; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_553 = 10'h229 == cpu_index ? cache_data_553 : _GEN_552; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_554 = 10'h22a == cpu_index ? cache_data_554 : _GEN_553; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_555 = 10'h22b == cpu_index ? cache_data_555 : _GEN_554; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_556 = 10'h22c == cpu_index ? cache_data_556 : _GEN_555; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_557 = 10'h22d == cpu_index ? cache_data_557 : _GEN_556; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_558 = 10'h22e == cpu_index ? cache_data_558 : _GEN_557; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_559 = 10'h22f == cpu_index ? cache_data_559 : _GEN_558; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_560 = 10'h230 == cpu_index ? cache_data_560 : _GEN_559; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_561 = 10'h231 == cpu_index ? cache_data_561 : _GEN_560; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_562 = 10'h232 == cpu_index ? cache_data_562 : _GEN_561; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_563 = 10'h233 == cpu_index ? cache_data_563 : _GEN_562; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_564 = 10'h234 == cpu_index ? cache_data_564 : _GEN_563; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_565 = 10'h235 == cpu_index ? cache_data_565 : _GEN_564; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_566 = 10'h236 == cpu_index ? cache_data_566 : _GEN_565; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_567 = 10'h237 == cpu_index ? cache_data_567 : _GEN_566; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_568 = 10'h238 == cpu_index ? cache_data_568 : _GEN_567; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_569 = 10'h239 == cpu_index ? cache_data_569 : _GEN_568; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_570 = 10'h23a == cpu_index ? cache_data_570 : _GEN_569; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_571 = 10'h23b == cpu_index ? cache_data_571 : _GEN_570; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_572 = 10'h23c == cpu_index ? cache_data_572 : _GEN_571; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_573 = 10'h23d == cpu_index ? cache_data_573 : _GEN_572; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_574 = 10'h23e == cpu_index ? cache_data_574 : _GEN_573; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_575 = 10'h23f == cpu_index ? cache_data_575 : _GEN_574; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_576 = 10'h240 == cpu_index ? cache_data_576 : _GEN_575; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_577 = 10'h241 == cpu_index ? cache_data_577 : _GEN_576; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_578 = 10'h242 == cpu_index ? cache_data_578 : _GEN_577; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_579 = 10'h243 == cpu_index ? cache_data_579 : _GEN_578; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_580 = 10'h244 == cpu_index ? cache_data_580 : _GEN_579; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_581 = 10'h245 == cpu_index ? cache_data_581 : _GEN_580; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_582 = 10'h246 == cpu_index ? cache_data_582 : _GEN_581; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_583 = 10'h247 == cpu_index ? cache_data_583 : _GEN_582; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_584 = 10'h248 == cpu_index ? cache_data_584 : _GEN_583; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_585 = 10'h249 == cpu_index ? cache_data_585 : _GEN_584; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_586 = 10'h24a == cpu_index ? cache_data_586 : _GEN_585; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_587 = 10'h24b == cpu_index ? cache_data_587 : _GEN_586; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_588 = 10'h24c == cpu_index ? cache_data_588 : _GEN_587; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_589 = 10'h24d == cpu_index ? cache_data_589 : _GEN_588; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_590 = 10'h24e == cpu_index ? cache_data_590 : _GEN_589; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_591 = 10'h24f == cpu_index ? cache_data_591 : _GEN_590; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_592 = 10'h250 == cpu_index ? cache_data_592 : _GEN_591; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_593 = 10'h251 == cpu_index ? cache_data_593 : _GEN_592; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_594 = 10'h252 == cpu_index ? cache_data_594 : _GEN_593; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_595 = 10'h253 == cpu_index ? cache_data_595 : _GEN_594; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_596 = 10'h254 == cpu_index ? cache_data_596 : _GEN_595; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_597 = 10'h255 == cpu_index ? cache_data_597 : _GEN_596; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_598 = 10'h256 == cpu_index ? cache_data_598 : _GEN_597; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_599 = 10'h257 == cpu_index ? cache_data_599 : _GEN_598; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_600 = 10'h258 == cpu_index ? cache_data_600 : _GEN_599; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_601 = 10'h259 == cpu_index ? cache_data_601 : _GEN_600; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_602 = 10'h25a == cpu_index ? cache_data_602 : _GEN_601; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_603 = 10'h25b == cpu_index ? cache_data_603 : _GEN_602; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_604 = 10'h25c == cpu_index ? cache_data_604 : _GEN_603; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_605 = 10'h25d == cpu_index ? cache_data_605 : _GEN_604; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_606 = 10'h25e == cpu_index ? cache_data_606 : _GEN_605; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_607 = 10'h25f == cpu_index ? cache_data_607 : _GEN_606; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_608 = 10'h260 == cpu_index ? cache_data_608 : _GEN_607; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_609 = 10'h261 == cpu_index ? cache_data_609 : _GEN_608; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_610 = 10'h262 == cpu_index ? cache_data_610 : _GEN_609; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_611 = 10'h263 == cpu_index ? cache_data_611 : _GEN_610; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_612 = 10'h264 == cpu_index ? cache_data_612 : _GEN_611; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_613 = 10'h265 == cpu_index ? cache_data_613 : _GEN_612; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_614 = 10'h266 == cpu_index ? cache_data_614 : _GEN_613; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_615 = 10'h267 == cpu_index ? cache_data_615 : _GEN_614; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_616 = 10'h268 == cpu_index ? cache_data_616 : _GEN_615; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_617 = 10'h269 == cpu_index ? cache_data_617 : _GEN_616; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_618 = 10'h26a == cpu_index ? cache_data_618 : _GEN_617; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_619 = 10'h26b == cpu_index ? cache_data_619 : _GEN_618; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_620 = 10'h26c == cpu_index ? cache_data_620 : _GEN_619; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_621 = 10'h26d == cpu_index ? cache_data_621 : _GEN_620; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_622 = 10'h26e == cpu_index ? cache_data_622 : _GEN_621; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_623 = 10'h26f == cpu_index ? cache_data_623 : _GEN_622; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_624 = 10'h270 == cpu_index ? cache_data_624 : _GEN_623; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_625 = 10'h271 == cpu_index ? cache_data_625 : _GEN_624; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_626 = 10'h272 == cpu_index ? cache_data_626 : _GEN_625; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_627 = 10'h273 == cpu_index ? cache_data_627 : _GEN_626; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_628 = 10'h274 == cpu_index ? cache_data_628 : _GEN_627; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_629 = 10'h275 == cpu_index ? cache_data_629 : _GEN_628; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_630 = 10'h276 == cpu_index ? cache_data_630 : _GEN_629; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_631 = 10'h277 == cpu_index ? cache_data_631 : _GEN_630; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_632 = 10'h278 == cpu_index ? cache_data_632 : _GEN_631; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_633 = 10'h279 == cpu_index ? cache_data_633 : _GEN_632; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_634 = 10'h27a == cpu_index ? cache_data_634 : _GEN_633; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_635 = 10'h27b == cpu_index ? cache_data_635 : _GEN_634; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_636 = 10'h27c == cpu_index ? cache_data_636 : _GEN_635; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_637 = 10'h27d == cpu_index ? cache_data_637 : _GEN_636; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_638 = 10'h27e == cpu_index ? cache_data_638 : _GEN_637; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_639 = 10'h27f == cpu_index ? cache_data_639 : _GEN_638; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_640 = 10'h280 == cpu_index ? cache_data_640 : _GEN_639; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_641 = 10'h281 == cpu_index ? cache_data_641 : _GEN_640; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_642 = 10'h282 == cpu_index ? cache_data_642 : _GEN_641; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_643 = 10'h283 == cpu_index ? cache_data_643 : _GEN_642; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_644 = 10'h284 == cpu_index ? cache_data_644 : _GEN_643; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_645 = 10'h285 == cpu_index ? cache_data_645 : _GEN_644; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_646 = 10'h286 == cpu_index ? cache_data_646 : _GEN_645; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_647 = 10'h287 == cpu_index ? cache_data_647 : _GEN_646; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_648 = 10'h288 == cpu_index ? cache_data_648 : _GEN_647; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_649 = 10'h289 == cpu_index ? cache_data_649 : _GEN_648; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_650 = 10'h28a == cpu_index ? cache_data_650 : _GEN_649; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_651 = 10'h28b == cpu_index ? cache_data_651 : _GEN_650; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_652 = 10'h28c == cpu_index ? cache_data_652 : _GEN_651; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_653 = 10'h28d == cpu_index ? cache_data_653 : _GEN_652; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_654 = 10'h28e == cpu_index ? cache_data_654 : _GEN_653; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_655 = 10'h28f == cpu_index ? cache_data_655 : _GEN_654; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_656 = 10'h290 == cpu_index ? cache_data_656 : _GEN_655; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_657 = 10'h291 == cpu_index ? cache_data_657 : _GEN_656; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_658 = 10'h292 == cpu_index ? cache_data_658 : _GEN_657; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_659 = 10'h293 == cpu_index ? cache_data_659 : _GEN_658; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_660 = 10'h294 == cpu_index ? cache_data_660 : _GEN_659; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_661 = 10'h295 == cpu_index ? cache_data_661 : _GEN_660; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_662 = 10'h296 == cpu_index ? cache_data_662 : _GEN_661; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_663 = 10'h297 == cpu_index ? cache_data_663 : _GEN_662; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_664 = 10'h298 == cpu_index ? cache_data_664 : _GEN_663; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_665 = 10'h299 == cpu_index ? cache_data_665 : _GEN_664; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_666 = 10'h29a == cpu_index ? cache_data_666 : _GEN_665; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_667 = 10'h29b == cpu_index ? cache_data_667 : _GEN_666; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_668 = 10'h29c == cpu_index ? cache_data_668 : _GEN_667; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_669 = 10'h29d == cpu_index ? cache_data_669 : _GEN_668; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_670 = 10'h29e == cpu_index ? cache_data_670 : _GEN_669; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_671 = 10'h29f == cpu_index ? cache_data_671 : _GEN_670; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_672 = 10'h2a0 == cpu_index ? cache_data_672 : _GEN_671; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_673 = 10'h2a1 == cpu_index ? cache_data_673 : _GEN_672; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_674 = 10'h2a2 == cpu_index ? cache_data_674 : _GEN_673; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_675 = 10'h2a3 == cpu_index ? cache_data_675 : _GEN_674; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_676 = 10'h2a4 == cpu_index ? cache_data_676 : _GEN_675; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_677 = 10'h2a5 == cpu_index ? cache_data_677 : _GEN_676; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_678 = 10'h2a6 == cpu_index ? cache_data_678 : _GEN_677; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_679 = 10'h2a7 == cpu_index ? cache_data_679 : _GEN_678; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_680 = 10'h2a8 == cpu_index ? cache_data_680 : _GEN_679; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_681 = 10'h2a9 == cpu_index ? cache_data_681 : _GEN_680; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_682 = 10'h2aa == cpu_index ? cache_data_682 : _GEN_681; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_683 = 10'h2ab == cpu_index ? cache_data_683 : _GEN_682; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_684 = 10'h2ac == cpu_index ? cache_data_684 : _GEN_683; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_685 = 10'h2ad == cpu_index ? cache_data_685 : _GEN_684; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_686 = 10'h2ae == cpu_index ? cache_data_686 : _GEN_685; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_687 = 10'h2af == cpu_index ? cache_data_687 : _GEN_686; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_688 = 10'h2b0 == cpu_index ? cache_data_688 : _GEN_687; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_689 = 10'h2b1 == cpu_index ? cache_data_689 : _GEN_688; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_690 = 10'h2b2 == cpu_index ? cache_data_690 : _GEN_689; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_691 = 10'h2b3 == cpu_index ? cache_data_691 : _GEN_690; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_692 = 10'h2b4 == cpu_index ? cache_data_692 : _GEN_691; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_693 = 10'h2b5 == cpu_index ? cache_data_693 : _GEN_692; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_694 = 10'h2b6 == cpu_index ? cache_data_694 : _GEN_693; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_695 = 10'h2b7 == cpu_index ? cache_data_695 : _GEN_694; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_696 = 10'h2b8 == cpu_index ? cache_data_696 : _GEN_695; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_697 = 10'h2b9 == cpu_index ? cache_data_697 : _GEN_696; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_698 = 10'h2ba == cpu_index ? cache_data_698 : _GEN_697; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_699 = 10'h2bb == cpu_index ? cache_data_699 : _GEN_698; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_700 = 10'h2bc == cpu_index ? cache_data_700 : _GEN_699; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_701 = 10'h2bd == cpu_index ? cache_data_701 : _GEN_700; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_702 = 10'h2be == cpu_index ? cache_data_702 : _GEN_701; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_703 = 10'h2bf == cpu_index ? cache_data_703 : _GEN_702; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_704 = 10'h2c0 == cpu_index ? cache_data_704 : _GEN_703; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_705 = 10'h2c1 == cpu_index ? cache_data_705 : _GEN_704; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_706 = 10'h2c2 == cpu_index ? cache_data_706 : _GEN_705; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_707 = 10'h2c3 == cpu_index ? cache_data_707 : _GEN_706; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_708 = 10'h2c4 == cpu_index ? cache_data_708 : _GEN_707; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_709 = 10'h2c5 == cpu_index ? cache_data_709 : _GEN_708; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_710 = 10'h2c6 == cpu_index ? cache_data_710 : _GEN_709; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_711 = 10'h2c7 == cpu_index ? cache_data_711 : _GEN_710; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_712 = 10'h2c8 == cpu_index ? cache_data_712 : _GEN_711; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_713 = 10'h2c9 == cpu_index ? cache_data_713 : _GEN_712; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_714 = 10'h2ca == cpu_index ? cache_data_714 : _GEN_713; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_715 = 10'h2cb == cpu_index ? cache_data_715 : _GEN_714; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_716 = 10'h2cc == cpu_index ? cache_data_716 : _GEN_715; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_717 = 10'h2cd == cpu_index ? cache_data_717 : _GEN_716; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_718 = 10'h2ce == cpu_index ? cache_data_718 : _GEN_717; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_719 = 10'h2cf == cpu_index ? cache_data_719 : _GEN_718; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_720 = 10'h2d0 == cpu_index ? cache_data_720 : _GEN_719; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_721 = 10'h2d1 == cpu_index ? cache_data_721 : _GEN_720; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_722 = 10'h2d2 == cpu_index ? cache_data_722 : _GEN_721; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_723 = 10'h2d3 == cpu_index ? cache_data_723 : _GEN_722; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_724 = 10'h2d4 == cpu_index ? cache_data_724 : _GEN_723; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_725 = 10'h2d5 == cpu_index ? cache_data_725 : _GEN_724; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_726 = 10'h2d6 == cpu_index ? cache_data_726 : _GEN_725; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_727 = 10'h2d7 == cpu_index ? cache_data_727 : _GEN_726; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_728 = 10'h2d8 == cpu_index ? cache_data_728 : _GEN_727; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_729 = 10'h2d9 == cpu_index ? cache_data_729 : _GEN_728; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_730 = 10'h2da == cpu_index ? cache_data_730 : _GEN_729; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_731 = 10'h2db == cpu_index ? cache_data_731 : _GEN_730; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_732 = 10'h2dc == cpu_index ? cache_data_732 : _GEN_731; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_733 = 10'h2dd == cpu_index ? cache_data_733 : _GEN_732; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_734 = 10'h2de == cpu_index ? cache_data_734 : _GEN_733; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_735 = 10'h2df == cpu_index ? cache_data_735 : _GEN_734; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_736 = 10'h2e0 == cpu_index ? cache_data_736 : _GEN_735; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_737 = 10'h2e1 == cpu_index ? cache_data_737 : _GEN_736; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_738 = 10'h2e2 == cpu_index ? cache_data_738 : _GEN_737; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_739 = 10'h2e3 == cpu_index ? cache_data_739 : _GEN_738; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_740 = 10'h2e4 == cpu_index ? cache_data_740 : _GEN_739; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_741 = 10'h2e5 == cpu_index ? cache_data_741 : _GEN_740; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_742 = 10'h2e6 == cpu_index ? cache_data_742 : _GEN_741; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_743 = 10'h2e7 == cpu_index ? cache_data_743 : _GEN_742; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_744 = 10'h2e8 == cpu_index ? cache_data_744 : _GEN_743; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_745 = 10'h2e9 == cpu_index ? cache_data_745 : _GEN_744; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_746 = 10'h2ea == cpu_index ? cache_data_746 : _GEN_745; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_747 = 10'h2eb == cpu_index ? cache_data_747 : _GEN_746; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_748 = 10'h2ec == cpu_index ? cache_data_748 : _GEN_747; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_749 = 10'h2ed == cpu_index ? cache_data_749 : _GEN_748; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_750 = 10'h2ee == cpu_index ? cache_data_750 : _GEN_749; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_751 = 10'h2ef == cpu_index ? cache_data_751 : _GEN_750; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_752 = 10'h2f0 == cpu_index ? cache_data_752 : _GEN_751; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_753 = 10'h2f1 == cpu_index ? cache_data_753 : _GEN_752; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_754 = 10'h2f2 == cpu_index ? cache_data_754 : _GEN_753; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_755 = 10'h2f3 == cpu_index ? cache_data_755 : _GEN_754; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_756 = 10'h2f4 == cpu_index ? cache_data_756 : _GEN_755; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_757 = 10'h2f5 == cpu_index ? cache_data_757 : _GEN_756; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_758 = 10'h2f6 == cpu_index ? cache_data_758 : _GEN_757; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_759 = 10'h2f7 == cpu_index ? cache_data_759 : _GEN_758; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_760 = 10'h2f8 == cpu_index ? cache_data_760 : _GEN_759; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_761 = 10'h2f9 == cpu_index ? cache_data_761 : _GEN_760; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_762 = 10'h2fa == cpu_index ? cache_data_762 : _GEN_761; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_763 = 10'h2fb == cpu_index ? cache_data_763 : _GEN_762; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_764 = 10'h2fc == cpu_index ? cache_data_764 : _GEN_763; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_765 = 10'h2fd == cpu_index ? cache_data_765 : _GEN_764; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_766 = 10'h2fe == cpu_index ? cache_data_766 : _GEN_765; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_767 = 10'h2ff == cpu_index ? cache_data_767 : _GEN_766; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_768 = 10'h300 == cpu_index ? cache_data_768 : _GEN_767; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_769 = 10'h301 == cpu_index ? cache_data_769 : _GEN_768; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_770 = 10'h302 == cpu_index ? cache_data_770 : _GEN_769; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_771 = 10'h303 == cpu_index ? cache_data_771 : _GEN_770; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_772 = 10'h304 == cpu_index ? cache_data_772 : _GEN_771; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_773 = 10'h305 == cpu_index ? cache_data_773 : _GEN_772; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_774 = 10'h306 == cpu_index ? cache_data_774 : _GEN_773; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_775 = 10'h307 == cpu_index ? cache_data_775 : _GEN_774; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_776 = 10'h308 == cpu_index ? cache_data_776 : _GEN_775; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_777 = 10'h309 == cpu_index ? cache_data_777 : _GEN_776; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_778 = 10'h30a == cpu_index ? cache_data_778 : _GEN_777; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_779 = 10'h30b == cpu_index ? cache_data_779 : _GEN_778; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_780 = 10'h30c == cpu_index ? cache_data_780 : _GEN_779; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_781 = 10'h30d == cpu_index ? cache_data_781 : _GEN_780; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_782 = 10'h30e == cpu_index ? cache_data_782 : _GEN_781; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_783 = 10'h30f == cpu_index ? cache_data_783 : _GEN_782; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_784 = 10'h310 == cpu_index ? cache_data_784 : _GEN_783; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_785 = 10'h311 == cpu_index ? cache_data_785 : _GEN_784; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_786 = 10'h312 == cpu_index ? cache_data_786 : _GEN_785; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_787 = 10'h313 == cpu_index ? cache_data_787 : _GEN_786; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_788 = 10'h314 == cpu_index ? cache_data_788 : _GEN_787; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_789 = 10'h315 == cpu_index ? cache_data_789 : _GEN_788; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_790 = 10'h316 == cpu_index ? cache_data_790 : _GEN_789; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_791 = 10'h317 == cpu_index ? cache_data_791 : _GEN_790; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_792 = 10'h318 == cpu_index ? cache_data_792 : _GEN_791; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_793 = 10'h319 == cpu_index ? cache_data_793 : _GEN_792; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_794 = 10'h31a == cpu_index ? cache_data_794 : _GEN_793; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_795 = 10'h31b == cpu_index ? cache_data_795 : _GEN_794; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_796 = 10'h31c == cpu_index ? cache_data_796 : _GEN_795; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_797 = 10'h31d == cpu_index ? cache_data_797 : _GEN_796; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_798 = 10'h31e == cpu_index ? cache_data_798 : _GEN_797; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_799 = 10'h31f == cpu_index ? cache_data_799 : _GEN_798; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_800 = 10'h320 == cpu_index ? cache_data_800 : _GEN_799; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_801 = 10'h321 == cpu_index ? cache_data_801 : _GEN_800; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_802 = 10'h322 == cpu_index ? cache_data_802 : _GEN_801; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_803 = 10'h323 == cpu_index ? cache_data_803 : _GEN_802; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_804 = 10'h324 == cpu_index ? cache_data_804 : _GEN_803; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_805 = 10'h325 == cpu_index ? cache_data_805 : _GEN_804; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_806 = 10'h326 == cpu_index ? cache_data_806 : _GEN_805; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_807 = 10'h327 == cpu_index ? cache_data_807 : _GEN_806; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_808 = 10'h328 == cpu_index ? cache_data_808 : _GEN_807; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_809 = 10'h329 == cpu_index ? cache_data_809 : _GEN_808; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_810 = 10'h32a == cpu_index ? cache_data_810 : _GEN_809; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_811 = 10'h32b == cpu_index ? cache_data_811 : _GEN_810; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_812 = 10'h32c == cpu_index ? cache_data_812 : _GEN_811; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_813 = 10'h32d == cpu_index ? cache_data_813 : _GEN_812; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_814 = 10'h32e == cpu_index ? cache_data_814 : _GEN_813; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_815 = 10'h32f == cpu_index ? cache_data_815 : _GEN_814; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_816 = 10'h330 == cpu_index ? cache_data_816 : _GEN_815; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_817 = 10'h331 == cpu_index ? cache_data_817 : _GEN_816; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_818 = 10'h332 == cpu_index ? cache_data_818 : _GEN_817; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_819 = 10'h333 == cpu_index ? cache_data_819 : _GEN_818; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_820 = 10'h334 == cpu_index ? cache_data_820 : _GEN_819; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_821 = 10'h335 == cpu_index ? cache_data_821 : _GEN_820; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_822 = 10'h336 == cpu_index ? cache_data_822 : _GEN_821; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_823 = 10'h337 == cpu_index ? cache_data_823 : _GEN_822; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_824 = 10'h338 == cpu_index ? cache_data_824 : _GEN_823; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_825 = 10'h339 == cpu_index ? cache_data_825 : _GEN_824; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_826 = 10'h33a == cpu_index ? cache_data_826 : _GEN_825; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_827 = 10'h33b == cpu_index ? cache_data_827 : _GEN_826; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_828 = 10'h33c == cpu_index ? cache_data_828 : _GEN_827; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_829 = 10'h33d == cpu_index ? cache_data_829 : _GEN_828; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_830 = 10'h33e == cpu_index ? cache_data_830 : _GEN_829; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_831 = 10'h33f == cpu_index ? cache_data_831 : _GEN_830; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_832 = 10'h340 == cpu_index ? cache_data_832 : _GEN_831; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_833 = 10'h341 == cpu_index ? cache_data_833 : _GEN_832; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_834 = 10'h342 == cpu_index ? cache_data_834 : _GEN_833; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_835 = 10'h343 == cpu_index ? cache_data_835 : _GEN_834; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_836 = 10'h344 == cpu_index ? cache_data_836 : _GEN_835; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_837 = 10'h345 == cpu_index ? cache_data_837 : _GEN_836; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_838 = 10'h346 == cpu_index ? cache_data_838 : _GEN_837; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_839 = 10'h347 == cpu_index ? cache_data_839 : _GEN_838; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_840 = 10'h348 == cpu_index ? cache_data_840 : _GEN_839; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_841 = 10'h349 == cpu_index ? cache_data_841 : _GEN_840; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_842 = 10'h34a == cpu_index ? cache_data_842 : _GEN_841; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_843 = 10'h34b == cpu_index ? cache_data_843 : _GEN_842; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_844 = 10'h34c == cpu_index ? cache_data_844 : _GEN_843; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_845 = 10'h34d == cpu_index ? cache_data_845 : _GEN_844; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_846 = 10'h34e == cpu_index ? cache_data_846 : _GEN_845; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_847 = 10'h34f == cpu_index ? cache_data_847 : _GEN_846; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_848 = 10'h350 == cpu_index ? cache_data_848 : _GEN_847; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_849 = 10'h351 == cpu_index ? cache_data_849 : _GEN_848; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_850 = 10'h352 == cpu_index ? cache_data_850 : _GEN_849; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_851 = 10'h353 == cpu_index ? cache_data_851 : _GEN_850; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_852 = 10'h354 == cpu_index ? cache_data_852 : _GEN_851; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_853 = 10'h355 == cpu_index ? cache_data_853 : _GEN_852; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_854 = 10'h356 == cpu_index ? cache_data_854 : _GEN_853; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_855 = 10'h357 == cpu_index ? cache_data_855 : _GEN_854; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_856 = 10'h358 == cpu_index ? cache_data_856 : _GEN_855; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_857 = 10'h359 == cpu_index ? cache_data_857 : _GEN_856; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_858 = 10'h35a == cpu_index ? cache_data_858 : _GEN_857; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_859 = 10'h35b == cpu_index ? cache_data_859 : _GEN_858; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_860 = 10'h35c == cpu_index ? cache_data_860 : _GEN_859; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_861 = 10'h35d == cpu_index ? cache_data_861 : _GEN_860; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_862 = 10'h35e == cpu_index ? cache_data_862 : _GEN_861; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_863 = 10'h35f == cpu_index ? cache_data_863 : _GEN_862; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_864 = 10'h360 == cpu_index ? cache_data_864 : _GEN_863; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_865 = 10'h361 == cpu_index ? cache_data_865 : _GEN_864; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_866 = 10'h362 == cpu_index ? cache_data_866 : _GEN_865; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_867 = 10'h363 == cpu_index ? cache_data_867 : _GEN_866; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_868 = 10'h364 == cpu_index ? cache_data_868 : _GEN_867; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_869 = 10'h365 == cpu_index ? cache_data_869 : _GEN_868; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_870 = 10'h366 == cpu_index ? cache_data_870 : _GEN_869; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_871 = 10'h367 == cpu_index ? cache_data_871 : _GEN_870; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_872 = 10'h368 == cpu_index ? cache_data_872 : _GEN_871; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_873 = 10'h369 == cpu_index ? cache_data_873 : _GEN_872; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_874 = 10'h36a == cpu_index ? cache_data_874 : _GEN_873; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_875 = 10'h36b == cpu_index ? cache_data_875 : _GEN_874; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_876 = 10'h36c == cpu_index ? cache_data_876 : _GEN_875; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_877 = 10'h36d == cpu_index ? cache_data_877 : _GEN_876; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_878 = 10'h36e == cpu_index ? cache_data_878 : _GEN_877; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_879 = 10'h36f == cpu_index ? cache_data_879 : _GEN_878; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_880 = 10'h370 == cpu_index ? cache_data_880 : _GEN_879; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_881 = 10'h371 == cpu_index ? cache_data_881 : _GEN_880; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_882 = 10'h372 == cpu_index ? cache_data_882 : _GEN_881; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_883 = 10'h373 == cpu_index ? cache_data_883 : _GEN_882; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_884 = 10'h374 == cpu_index ? cache_data_884 : _GEN_883; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_885 = 10'h375 == cpu_index ? cache_data_885 : _GEN_884; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_886 = 10'h376 == cpu_index ? cache_data_886 : _GEN_885; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_887 = 10'h377 == cpu_index ? cache_data_887 : _GEN_886; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_888 = 10'h378 == cpu_index ? cache_data_888 : _GEN_887; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_889 = 10'h379 == cpu_index ? cache_data_889 : _GEN_888; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_890 = 10'h37a == cpu_index ? cache_data_890 : _GEN_889; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_891 = 10'h37b == cpu_index ? cache_data_891 : _GEN_890; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_892 = 10'h37c == cpu_index ? cache_data_892 : _GEN_891; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_893 = 10'h37d == cpu_index ? cache_data_893 : _GEN_892; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_894 = 10'h37e == cpu_index ? cache_data_894 : _GEN_893; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_895 = 10'h37f == cpu_index ? cache_data_895 : _GEN_894; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_896 = 10'h380 == cpu_index ? cache_data_896 : _GEN_895; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_897 = 10'h381 == cpu_index ? cache_data_897 : _GEN_896; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_898 = 10'h382 == cpu_index ? cache_data_898 : _GEN_897; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_899 = 10'h383 == cpu_index ? cache_data_899 : _GEN_898; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_900 = 10'h384 == cpu_index ? cache_data_900 : _GEN_899; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_901 = 10'h385 == cpu_index ? cache_data_901 : _GEN_900; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_902 = 10'h386 == cpu_index ? cache_data_902 : _GEN_901; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_903 = 10'h387 == cpu_index ? cache_data_903 : _GEN_902; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_904 = 10'h388 == cpu_index ? cache_data_904 : _GEN_903; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_905 = 10'h389 == cpu_index ? cache_data_905 : _GEN_904; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_906 = 10'h38a == cpu_index ? cache_data_906 : _GEN_905; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_907 = 10'h38b == cpu_index ? cache_data_907 : _GEN_906; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_908 = 10'h38c == cpu_index ? cache_data_908 : _GEN_907; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_909 = 10'h38d == cpu_index ? cache_data_909 : _GEN_908; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_910 = 10'h38e == cpu_index ? cache_data_910 : _GEN_909; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_911 = 10'h38f == cpu_index ? cache_data_911 : _GEN_910; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_912 = 10'h390 == cpu_index ? cache_data_912 : _GEN_911; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_913 = 10'h391 == cpu_index ? cache_data_913 : _GEN_912; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_914 = 10'h392 == cpu_index ? cache_data_914 : _GEN_913; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_915 = 10'h393 == cpu_index ? cache_data_915 : _GEN_914; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_916 = 10'h394 == cpu_index ? cache_data_916 : _GEN_915; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_917 = 10'h395 == cpu_index ? cache_data_917 : _GEN_916; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_918 = 10'h396 == cpu_index ? cache_data_918 : _GEN_917; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_919 = 10'h397 == cpu_index ? cache_data_919 : _GEN_918; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_920 = 10'h398 == cpu_index ? cache_data_920 : _GEN_919; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_921 = 10'h399 == cpu_index ? cache_data_921 : _GEN_920; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_922 = 10'h39a == cpu_index ? cache_data_922 : _GEN_921; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_923 = 10'h39b == cpu_index ? cache_data_923 : _GEN_922; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_924 = 10'h39c == cpu_index ? cache_data_924 : _GEN_923; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_925 = 10'h39d == cpu_index ? cache_data_925 : _GEN_924; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_926 = 10'h39e == cpu_index ? cache_data_926 : _GEN_925; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_927 = 10'h39f == cpu_index ? cache_data_927 : _GEN_926; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_928 = 10'h3a0 == cpu_index ? cache_data_928 : _GEN_927; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_929 = 10'h3a1 == cpu_index ? cache_data_929 : _GEN_928; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_930 = 10'h3a2 == cpu_index ? cache_data_930 : _GEN_929; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_931 = 10'h3a3 == cpu_index ? cache_data_931 : _GEN_930; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_932 = 10'h3a4 == cpu_index ? cache_data_932 : _GEN_931; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_933 = 10'h3a5 == cpu_index ? cache_data_933 : _GEN_932; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_934 = 10'h3a6 == cpu_index ? cache_data_934 : _GEN_933; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_935 = 10'h3a7 == cpu_index ? cache_data_935 : _GEN_934; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_936 = 10'h3a8 == cpu_index ? cache_data_936 : _GEN_935; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_937 = 10'h3a9 == cpu_index ? cache_data_937 : _GEN_936; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_938 = 10'h3aa == cpu_index ? cache_data_938 : _GEN_937; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_939 = 10'h3ab == cpu_index ? cache_data_939 : _GEN_938; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_940 = 10'h3ac == cpu_index ? cache_data_940 : _GEN_939; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_941 = 10'h3ad == cpu_index ? cache_data_941 : _GEN_940; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_942 = 10'h3ae == cpu_index ? cache_data_942 : _GEN_941; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_943 = 10'h3af == cpu_index ? cache_data_943 : _GEN_942; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_944 = 10'h3b0 == cpu_index ? cache_data_944 : _GEN_943; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_945 = 10'h3b1 == cpu_index ? cache_data_945 : _GEN_944; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_946 = 10'h3b2 == cpu_index ? cache_data_946 : _GEN_945; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_947 = 10'h3b3 == cpu_index ? cache_data_947 : _GEN_946; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_948 = 10'h3b4 == cpu_index ? cache_data_948 : _GEN_947; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_949 = 10'h3b5 == cpu_index ? cache_data_949 : _GEN_948; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_950 = 10'h3b6 == cpu_index ? cache_data_950 : _GEN_949; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_951 = 10'h3b7 == cpu_index ? cache_data_951 : _GEN_950; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_952 = 10'h3b8 == cpu_index ? cache_data_952 : _GEN_951; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_953 = 10'h3b9 == cpu_index ? cache_data_953 : _GEN_952; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_954 = 10'h3ba == cpu_index ? cache_data_954 : _GEN_953; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_955 = 10'h3bb == cpu_index ? cache_data_955 : _GEN_954; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_956 = 10'h3bc == cpu_index ? cache_data_956 : _GEN_955; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_957 = 10'h3bd == cpu_index ? cache_data_957 : _GEN_956; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_958 = 10'h3be == cpu_index ? cache_data_958 : _GEN_957; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_959 = 10'h3bf == cpu_index ? cache_data_959 : _GEN_958; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_960 = 10'h3c0 == cpu_index ? cache_data_960 : _GEN_959; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_961 = 10'h3c1 == cpu_index ? cache_data_961 : _GEN_960; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_962 = 10'h3c2 == cpu_index ? cache_data_962 : _GEN_961; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_963 = 10'h3c3 == cpu_index ? cache_data_963 : _GEN_962; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_964 = 10'h3c4 == cpu_index ? cache_data_964 : _GEN_963; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_965 = 10'h3c5 == cpu_index ? cache_data_965 : _GEN_964; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_966 = 10'h3c6 == cpu_index ? cache_data_966 : _GEN_965; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_967 = 10'h3c7 == cpu_index ? cache_data_967 : _GEN_966; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_968 = 10'h3c8 == cpu_index ? cache_data_968 : _GEN_967; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_969 = 10'h3c9 == cpu_index ? cache_data_969 : _GEN_968; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_970 = 10'h3ca == cpu_index ? cache_data_970 : _GEN_969; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_971 = 10'h3cb == cpu_index ? cache_data_971 : _GEN_970; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_972 = 10'h3cc == cpu_index ? cache_data_972 : _GEN_971; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_973 = 10'h3cd == cpu_index ? cache_data_973 : _GEN_972; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_974 = 10'h3ce == cpu_index ? cache_data_974 : _GEN_973; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_975 = 10'h3cf == cpu_index ? cache_data_975 : _GEN_974; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_976 = 10'h3d0 == cpu_index ? cache_data_976 : _GEN_975; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_977 = 10'h3d1 == cpu_index ? cache_data_977 : _GEN_976; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_978 = 10'h3d2 == cpu_index ? cache_data_978 : _GEN_977; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_979 = 10'h3d3 == cpu_index ? cache_data_979 : _GEN_978; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_980 = 10'h3d4 == cpu_index ? cache_data_980 : _GEN_979; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_981 = 10'h3d5 == cpu_index ? cache_data_981 : _GEN_980; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_982 = 10'h3d6 == cpu_index ? cache_data_982 : _GEN_981; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_983 = 10'h3d7 == cpu_index ? cache_data_983 : _GEN_982; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_984 = 10'h3d8 == cpu_index ? cache_data_984 : _GEN_983; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_985 = 10'h3d9 == cpu_index ? cache_data_985 : _GEN_984; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_986 = 10'h3da == cpu_index ? cache_data_986 : _GEN_985; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_987 = 10'h3db == cpu_index ? cache_data_987 : _GEN_986; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_988 = 10'h3dc == cpu_index ? cache_data_988 : _GEN_987; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_989 = 10'h3dd == cpu_index ? cache_data_989 : _GEN_988; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_990 = 10'h3de == cpu_index ? cache_data_990 : _GEN_989; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_991 = 10'h3df == cpu_index ? cache_data_991 : _GEN_990; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_992 = 10'h3e0 == cpu_index ? cache_data_992 : _GEN_991; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_993 = 10'h3e1 == cpu_index ? cache_data_993 : _GEN_992; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_994 = 10'h3e2 == cpu_index ? cache_data_994 : _GEN_993; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_995 = 10'h3e3 == cpu_index ? cache_data_995 : _GEN_994; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_996 = 10'h3e4 == cpu_index ? cache_data_996 : _GEN_995; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_997 = 10'h3e5 == cpu_index ? cache_data_997 : _GEN_996; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_998 = 10'h3e6 == cpu_index ? cache_data_998 : _GEN_997; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_999 = 10'h3e7 == cpu_index ? cache_data_999 : _GEN_998; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1000 = 10'h3e8 == cpu_index ? cache_data_1000 : _GEN_999; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1001 = 10'h3e9 == cpu_index ? cache_data_1001 : _GEN_1000; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1002 = 10'h3ea == cpu_index ? cache_data_1002 : _GEN_1001; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1003 = 10'h3eb == cpu_index ? cache_data_1003 : _GEN_1002; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1004 = 10'h3ec == cpu_index ? cache_data_1004 : _GEN_1003; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1005 = 10'h3ed == cpu_index ? cache_data_1005 : _GEN_1004; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1006 = 10'h3ee == cpu_index ? cache_data_1006 : _GEN_1005; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1007 = 10'h3ef == cpu_index ? cache_data_1007 : _GEN_1006; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1008 = 10'h3f0 == cpu_index ? cache_data_1008 : _GEN_1007; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1009 = 10'h3f1 == cpu_index ? cache_data_1009 : _GEN_1008; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1010 = 10'h3f2 == cpu_index ? cache_data_1010 : _GEN_1009; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1011 = 10'h3f3 == cpu_index ? cache_data_1011 : _GEN_1010; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1012 = 10'h3f4 == cpu_index ? cache_data_1012 : _GEN_1011; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1013 = 10'h3f5 == cpu_index ? cache_data_1013 : _GEN_1012; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1014 = 10'h3f6 == cpu_index ? cache_data_1014 : _GEN_1013; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1015 = 10'h3f7 == cpu_index ? cache_data_1015 : _GEN_1014; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1016 = 10'h3f8 == cpu_index ? cache_data_1016 : _GEN_1015; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1017 = 10'h3f9 == cpu_index ? cache_data_1017 : _GEN_1016; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1018 = 10'h3fa == cpu_index ? cache_data_1018 : _GEN_1017; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1019 = 10'h3fb == cpu_index ? cache_data_1019 : _GEN_1018; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1020 = 10'h3fc == cpu_index ? cache_data_1020 : _GEN_1019; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1021 = 10'h3fd == cpu_index ? cache_data_1021 : _GEN_1020; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1022 = 10'h3fe == cpu_index ? cache_data_1022 : _GEN_1021; // @[icache.scala 48:{37,37}]
  wire [184:0] _GEN_1023 = 10'h3ff == cpu_index ? cache_data_1023 : _GEN_1022; // @[icache.scala 48:{37,37}]
  wire  way0_hit = _GEN_1023[184] & _GEN_1023[182:128] == cpu_tag; // @[icache.scala 48:52]
  wire [9:0] _way1_hit_T_1 = cpu_index + 10'h1; // @[icache.scala 49:37]
  wire [184:0] _GEN_1025 = 10'h1 == _way1_hit_T_1 ? cache_data_1 : cache_data_0; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1026 = 10'h2 == _way1_hit_T_1 ? cache_data_2 : _GEN_1025; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1027 = 10'h3 == _way1_hit_T_1 ? cache_data_3 : _GEN_1026; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1028 = 10'h4 == _way1_hit_T_1 ? cache_data_4 : _GEN_1027; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1029 = 10'h5 == _way1_hit_T_1 ? cache_data_5 : _GEN_1028; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1030 = 10'h6 == _way1_hit_T_1 ? cache_data_6 : _GEN_1029; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1031 = 10'h7 == _way1_hit_T_1 ? cache_data_7 : _GEN_1030; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1032 = 10'h8 == _way1_hit_T_1 ? cache_data_8 : _GEN_1031; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1033 = 10'h9 == _way1_hit_T_1 ? cache_data_9 : _GEN_1032; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1034 = 10'ha == _way1_hit_T_1 ? cache_data_10 : _GEN_1033; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1035 = 10'hb == _way1_hit_T_1 ? cache_data_11 : _GEN_1034; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1036 = 10'hc == _way1_hit_T_1 ? cache_data_12 : _GEN_1035; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1037 = 10'hd == _way1_hit_T_1 ? cache_data_13 : _GEN_1036; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1038 = 10'he == _way1_hit_T_1 ? cache_data_14 : _GEN_1037; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1039 = 10'hf == _way1_hit_T_1 ? cache_data_15 : _GEN_1038; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1040 = 10'h10 == _way1_hit_T_1 ? cache_data_16 : _GEN_1039; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1041 = 10'h11 == _way1_hit_T_1 ? cache_data_17 : _GEN_1040; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1042 = 10'h12 == _way1_hit_T_1 ? cache_data_18 : _GEN_1041; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1043 = 10'h13 == _way1_hit_T_1 ? cache_data_19 : _GEN_1042; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1044 = 10'h14 == _way1_hit_T_1 ? cache_data_20 : _GEN_1043; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1045 = 10'h15 == _way1_hit_T_1 ? cache_data_21 : _GEN_1044; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1046 = 10'h16 == _way1_hit_T_1 ? cache_data_22 : _GEN_1045; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1047 = 10'h17 == _way1_hit_T_1 ? cache_data_23 : _GEN_1046; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1048 = 10'h18 == _way1_hit_T_1 ? cache_data_24 : _GEN_1047; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1049 = 10'h19 == _way1_hit_T_1 ? cache_data_25 : _GEN_1048; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1050 = 10'h1a == _way1_hit_T_1 ? cache_data_26 : _GEN_1049; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1051 = 10'h1b == _way1_hit_T_1 ? cache_data_27 : _GEN_1050; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1052 = 10'h1c == _way1_hit_T_1 ? cache_data_28 : _GEN_1051; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1053 = 10'h1d == _way1_hit_T_1 ? cache_data_29 : _GEN_1052; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1054 = 10'h1e == _way1_hit_T_1 ? cache_data_30 : _GEN_1053; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1055 = 10'h1f == _way1_hit_T_1 ? cache_data_31 : _GEN_1054; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1056 = 10'h20 == _way1_hit_T_1 ? cache_data_32 : _GEN_1055; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1057 = 10'h21 == _way1_hit_T_1 ? cache_data_33 : _GEN_1056; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1058 = 10'h22 == _way1_hit_T_1 ? cache_data_34 : _GEN_1057; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1059 = 10'h23 == _way1_hit_T_1 ? cache_data_35 : _GEN_1058; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1060 = 10'h24 == _way1_hit_T_1 ? cache_data_36 : _GEN_1059; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1061 = 10'h25 == _way1_hit_T_1 ? cache_data_37 : _GEN_1060; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1062 = 10'h26 == _way1_hit_T_1 ? cache_data_38 : _GEN_1061; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1063 = 10'h27 == _way1_hit_T_1 ? cache_data_39 : _GEN_1062; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1064 = 10'h28 == _way1_hit_T_1 ? cache_data_40 : _GEN_1063; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1065 = 10'h29 == _way1_hit_T_1 ? cache_data_41 : _GEN_1064; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1066 = 10'h2a == _way1_hit_T_1 ? cache_data_42 : _GEN_1065; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1067 = 10'h2b == _way1_hit_T_1 ? cache_data_43 : _GEN_1066; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1068 = 10'h2c == _way1_hit_T_1 ? cache_data_44 : _GEN_1067; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1069 = 10'h2d == _way1_hit_T_1 ? cache_data_45 : _GEN_1068; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1070 = 10'h2e == _way1_hit_T_1 ? cache_data_46 : _GEN_1069; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1071 = 10'h2f == _way1_hit_T_1 ? cache_data_47 : _GEN_1070; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1072 = 10'h30 == _way1_hit_T_1 ? cache_data_48 : _GEN_1071; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1073 = 10'h31 == _way1_hit_T_1 ? cache_data_49 : _GEN_1072; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1074 = 10'h32 == _way1_hit_T_1 ? cache_data_50 : _GEN_1073; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1075 = 10'h33 == _way1_hit_T_1 ? cache_data_51 : _GEN_1074; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1076 = 10'h34 == _way1_hit_T_1 ? cache_data_52 : _GEN_1075; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1077 = 10'h35 == _way1_hit_T_1 ? cache_data_53 : _GEN_1076; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1078 = 10'h36 == _way1_hit_T_1 ? cache_data_54 : _GEN_1077; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1079 = 10'h37 == _way1_hit_T_1 ? cache_data_55 : _GEN_1078; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1080 = 10'h38 == _way1_hit_T_1 ? cache_data_56 : _GEN_1079; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1081 = 10'h39 == _way1_hit_T_1 ? cache_data_57 : _GEN_1080; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1082 = 10'h3a == _way1_hit_T_1 ? cache_data_58 : _GEN_1081; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1083 = 10'h3b == _way1_hit_T_1 ? cache_data_59 : _GEN_1082; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1084 = 10'h3c == _way1_hit_T_1 ? cache_data_60 : _GEN_1083; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1085 = 10'h3d == _way1_hit_T_1 ? cache_data_61 : _GEN_1084; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1086 = 10'h3e == _way1_hit_T_1 ? cache_data_62 : _GEN_1085; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1087 = 10'h3f == _way1_hit_T_1 ? cache_data_63 : _GEN_1086; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1088 = 10'h40 == _way1_hit_T_1 ? cache_data_64 : _GEN_1087; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1089 = 10'h41 == _way1_hit_T_1 ? cache_data_65 : _GEN_1088; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1090 = 10'h42 == _way1_hit_T_1 ? cache_data_66 : _GEN_1089; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1091 = 10'h43 == _way1_hit_T_1 ? cache_data_67 : _GEN_1090; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1092 = 10'h44 == _way1_hit_T_1 ? cache_data_68 : _GEN_1091; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1093 = 10'h45 == _way1_hit_T_1 ? cache_data_69 : _GEN_1092; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1094 = 10'h46 == _way1_hit_T_1 ? cache_data_70 : _GEN_1093; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1095 = 10'h47 == _way1_hit_T_1 ? cache_data_71 : _GEN_1094; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1096 = 10'h48 == _way1_hit_T_1 ? cache_data_72 : _GEN_1095; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1097 = 10'h49 == _way1_hit_T_1 ? cache_data_73 : _GEN_1096; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1098 = 10'h4a == _way1_hit_T_1 ? cache_data_74 : _GEN_1097; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1099 = 10'h4b == _way1_hit_T_1 ? cache_data_75 : _GEN_1098; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1100 = 10'h4c == _way1_hit_T_1 ? cache_data_76 : _GEN_1099; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1101 = 10'h4d == _way1_hit_T_1 ? cache_data_77 : _GEN_1100; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1102 = 10'h4e == _way1_hit_T_1 ? cache_data_78 : _GEN_1101; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1103 = 10'h4f == _way1_hit_T_1 ? cache_data_79 : _GEN_1102; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1104 = 10'h50 == _way1_hit_T_1 ? cache_data_80 : _GEN_1103; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1105 = 10'h51 == _way1_hit_T_1 ? cache_data_81 : _GEN_1104; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1106 = 10'h52 == _way1_hit_T_1 ? cache_data_82 : _GEN_1105; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1107 = 10'h53 == _way1_hit_T_1 ? cache_data_83 : _GEN_1106; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1108 = 10'h54 == _way1_hit_T_1 ? cache_data_84 : _GEN_1107; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1109 = 10'h55 == _way1_hit_T_1 ? cache_data_85 : _GEN_1108; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1110 = 10'h56 == _way1_hit_T_1 ? cache_data_86 : _GEN_1109; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1111 = 10'h57 == _way1_hit_T_1 ? cache_data_87 : _GEN_1110; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1112 = 10'h58 == _way1_hit_T_1 ? cache_data_88 : _GEN_1111; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1113 = 10'h59 == _way1_hit_T_1 ? cache_data_89 : _GEN_1112; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1114 = 10'h5a == _way1_hit_T_1 ? cache_data_90 : _GEN_1113; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1115 = 10'h5b == _way1_hit_T_1 ? cache_data_91 : _GEN_1114; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1116 = 10'h5c == _way1_hit_T_1 ? cache_data_92 : _GEN_1115; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1117 = 10'h5d == _way1_hit_T_1 ? cache_data_93 : _GEN_1116; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1118 = 10'h5e == _way1_hit_T_1 ? cache_data_94 : _GEN_1117; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1119 = 10'h5f == _way1_hit_T_1 ? cache_data_95 : _GEN_1118; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1120 = 10'h60 == _way1_hit_T_1 ? cache_data_96 : _GEN_1119; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1121 = 10'h61 == _way1_hit_T_1 ? cache_data_97 : _GEN_1120; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1122 = 10'h62 == _way1_hit_T_1 ? cache_data_98 : _GEN_1121; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1123 = 10'h63 == _way1_hit_T_1 ? cache_data_99 : _GEN_1122; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1124 = 10'h64 == _way1_hit_T_1 ? cache_data_100 : _GEN_1123; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1125 = 10'h65 == _way1_hit_T_1 ? cache_data_101 : _GEN_1124; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1126 = 10'h66 == _way1_hit_T_1 ? cache_data_102 : _GEN_1125; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1127 = 10'h67 == _way1_hit_T_1 ? cache_data_103 : _GEN_1126; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1128 = 10'h68 == _way1_hit_T_1 ? cache_data_104 : _GEN_1127; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1129 = 10'h69 == _way1_hit_T_1 ? cache_data_105 : _GEN_1128; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1130 = 10'h6a == _way1_hit_T_1 ? cache_data_106 : _GEN_1129; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1131 = 10'h6b == _way1_hit_T_1 ? cache_data_107 : _GEN_1130; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1132 = 10'h6c == _way1_hit_T_1 ? cache_data_108 : _GEN_1131; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1133 = 10'h6d == _way1_hit_T_1 ? cache_data_109 : _GEN_1132; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1134 = 10'h6e == _way1_hit_T_1 ? cache_data_110 : _GEN_1133; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1135 = 10'h6f == _way1_hit_T_1 ? cache_data_111 : _GEN_1134; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1136 = 10'h70 == _way1_hit_T_1 ? cache_data_112 : _GEN_1135; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1137 = 10'h71 == _way1_hit_T_1 ? cache_data_113 : _GEN_1136; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1138 = 10'h72 == _way1_hit_T_1 ? cache_data_114 : _GEN_1137; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1139 = 10'h73 == _way1_hit_T_1 ? cache_data_115 : _GEN_1138; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1140 = 10'h74 == _way1_hit_T_1 ? cache_data_116 : _GEN_1139; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1141 = 10'h75 == _way1_hit_T_1 ? cache_data_117 : _GEN_1140; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1142 = 10'h76 == _way1_hit_T_1 ? cache_data_118 : _GEN_1141; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1143 = 10'h77 == _way1_hit_T_1 ? cache_data_119 : _GEN_1142; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1144 = 10'h78 == _way1_hit_T_1 ? cache_data_120 : _GEN_1143; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1145 = 10'h79 == _way1_hit_T_1 ? cache_data_121 : _GEN_1144; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1146 = 10'h7a == _way1_hit_T_1 ? cache_data_122 : _GEN_1145; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1147 = 10'h7b == _way1_hit_T_1 ? cache_data_123 : _GEN_1146; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1148 = 10'h7c == _way1_hit_T_1 ? cache_data_124 : _GEN_1147; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1149 = 10'h7d == _way1_hit_T_1 ? cache_data_125 : _GEN_1148; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1150 = 10'h7e == _way1_hit_T_1 ? cache_data_126 : _GEN_1149; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1151 = 10'h7f == _way1_hit_T_1 ? cache_data_127 : _GEN_1150; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1152 = 10'h80 == _way1_hit_T_1 ? cache_data_128 : _GEN_1151; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1153 = 10'h81 == _way1_hit_T_1 ? cache_data_129 : _GEN_1152; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1154 = 10'h82 == _way1_hit_T_1 ? cache_data_130 : _GEN_1153; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1155 = 10'h83 == _way1_hit_T_1 ? cache_data_131 : _GEN_1154; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1156 = 10'h84 == _way1_hit_T_1 ? cache_data_132 : _GEN_1155; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1157 = 10'h85 == _way1_hit_T_1 ? cache_data_133 : _GEN_1156; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1158 = 10'h86 == _way1_hit_T_1 ? cache_data_134 : _GEN_1157; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1159 = 10'h87 == _way1_hit_T_1 ? cache_data_135 : _GEN_1158; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1160 = 10'h88 == _way1_hit_T_1 ? cache_data_136 : _GEN_1159; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1161 = 10'h89 == _way1_hit_T_1 ? cache_data_137 : _GEN_1160; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1162 = 10'h8a == _way1_hit_T_1 ? cache_data_138 : _GEN_1161; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1163 = 10'h8b == _way1_hit_T_1 ? cache_data_139 : _GEN_1162; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1164 = 10'h8c == _way1_hit_T_1 ? cache_data_140 : _GEN_1163; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1165 = 10'h8d == _way1_hit_T_1 ? cache_data_141 : _GEN_1164; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1166 = 10'h8e == _way1_hit_T_1 ? cache_data_142 : _GEN_1165; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1167 = 10'h8f == _way1_hit_T_1 ? cache_data_143 : _GEN_1166; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1168 = 10'h90 == _way1_hit_T_1 ? cache_data_144 : _GEN_1167; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1169 = 10'h91 == _way1_hit_T_1 ? cache_data_145 : _GEN_1168; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1170 = 10'h92 == _way1_hit_T_1 ? cache_data_146 : _GEN_1169; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1171 = 10'h93 == _way1_hit_T_1 ? cache_data_147 : _GEN_1170; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1172 = 10'h94 == _way1_hit_T_1 ? cache_data_148 : _GEN_1171; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1173 = 10'h95 == _way1_hit_T_1 ? cache_data_149 : _GEN_1172; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1174 = 10'h96 == _way1_hit_T_1 ? cache_data_150 : _GEN_1173; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1175 = 10'h97 == _way1_hit_T_1 ? cache_data_151 : _GEN_1174; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1176 = 10'h98 == _way1_hit_T_1 ? cache_data_152 : _GEN_1175; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1177 = 10'h99 == _way1_hit_T_1 ? cache_data_153 : _GEN_1176; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1178 = 10'h9a == _way1_hit_T_1 ? cache_data_154 : _GEN_1177; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1179 = 10'h9b == _way1_hit_T_1 ? cache_data_155 : _GEN_1178; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1180 = 10'h9c == _way1_hit_T_1 ? cache_data_156 : _GEN_1179; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1181 = 10'h9d == _way1_hit_T_1 ? cache_data_157 : _GEN_1180; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1182 = 10'h9e == _way1_hit_T_1 ? cache_data_158 : _GEN_1181; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1183 = 10'h9f == _way1_hit_T_1 ? cache_data_159 : _GEN_1182; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1184 = 10'ha0 == _way1_hit_T_1 ? cache_data_160 : _GEN_1183; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1185 = 10'ha1 == _way1_hit_T_1 ? cache_data_161 : _GEN_1184; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1186 = 10'ha2 == _way1_hit_T_1 ? cache_data_162 : _GEN_1185; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1187 = 10'ha3 == _way1_hit_T_1 ? cache_data_163 : _GEN_1186; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1188 = 10'ha4 == _way1_hit_T_1 ? cache_data_164 : _GEN_1187; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1189 = 10'ha5 == _way1_hit_T_1 ? cache_data_165 : _GEN_1188; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1190 = 10'ha6 == _way1_hit_T_1 ? cache_data_166 : _GEN_1189; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1191 = 10'ha7 == _way1_hit_T_1 ? cache_data_167 : _GEN_1190; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1192 = 10'ha8 == _way1_hit_T_1 ? cache_data_168 : _GEN_1191; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1193 = 10'ha9 == _way1_hit_T_1 ? cache_data_169 : _GEN_1192; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1194 = 10'haa == _way1_hit_T_1 ? cache_data_170 : _GEN_1193; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1195 = 10'hab == _way1_hit_T_1 ? cache_data_171 : _GEN_1194; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1196 = 10'hac == _way1_hit_T_1 ? cache_data_172 : _GEN_1195; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1197 = 10'had == _way1_hit_T_1 ? cache_data_173 : _GEN_1196; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1198 = 10'hae == _way1_hit_T_1 ? cache_data_174 : _GEN_1197; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1199 = 10'haf == _way1_hit_T_1 ? cache_data_175 : _GEN_1198; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1200 = 10'hb0 == _way1_hit_T_1 ? cache_data_176 : _GEN_1199; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1201 = 10'hb1 == _way1_hit_T_1 ? cache_data_177 : _GEN_1200; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1202 = 10'hb2 == _way1_hit_T_1 ? cache_data_178 : _GEN_1201; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1203 = 10'hb3 == _way1_hit_T_1 ? cache_data_179 : _GEN_1202; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1204 = 10'hb4 == _way1_hit_T_1 ? cache_data_180 : _GEN_1203; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1205 = 10'hb5 == _way1_hit_T_1 ? cache_data_181 : _GEN_1204; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1206 = 10'hb6 == _way1_hit_T_1 ? cache_data_182 : _GEN_1205; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1207 = 10'hb7 == _way1_hit_T_1 ? cache_data_183 : _GEN_1206; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1208 = 10'hb8 == _way1_hit_T_1 ? cache_data_184 : _GEN_1207; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1209 = 10'hb9 == _way1_hit_T_1 ? cache_data_185 : _GEN_1208; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1210 = 10'hba == _way1_hit_T_1 ? cache_data_186 : _GEN_1209; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1211 = 10'hbb == _way1_hit_T_1 ? cache_data_187 : _GEN_1210; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1212 = 10'hbc == _way1_hit_T_1 ? cache_data_188 : _GEN_1211; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1213 = 10'hbd == _way1_hit_T_1 ? cache_data_189 : _GEN_1212; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1214 = 10'hbe == _way1_hit_T_1 ? cache_data_190 : _GEN_1213; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1215 = 10'hbf == _way1_hit_T_1 ? cache_data_191 : _GEN_1214; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1216 = 10'hc0 == _way1_hit_T_1 ? cache_data_192 : _GEN_1215; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1217 = 10'hc1 == _way1_hit_T_1 ? cache_data_193 : _GEN_1216; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1218 = 10'hc2 == _way1_hit_T_1 ? cache_data_194 : _GEN_1217; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1219 = 10'hc3 == _way1_hit_T_1 ? cache_data_195 : _GEN_1218; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1220 = 10'hc4 == _way1_hit_T_1 ? cache_data_196 : _GEN_1219; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1221 = 10'hc5 == _way1_hit_T_1 ? cache_data_197 : _GEN_1220; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1222 = 10'hc6 == _way1_hit_T_1 ? cache_data_198 : _GEN_1221; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1223 = 10'hc7 == _way1_hit_T_1 ? cache_data_199 : _GEN_1222; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1224 = 10'hc8 == _way1_hit_T_1 ? cache_data_200 : _GEN_1223; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1225 = 10'hc9 == _way1_hit_T_1 ? cache_data_201 : _GEN_1224; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1226 = 10'hca == _way1_hit_T_1 ? cache_data_202 : _GEN_1225; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1227 = 10'hcb == _way1_hit_T_1 ? cache_data_203 : _GEN_1226; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1228 = 10'hcc == _way1_hit_T_1 ? cache_data_204 : _GEN_1227; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1229 = 10'hcd == _way1_hit_T_1 ? cache_data_205 : _GEN_1228; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1230 = 10'hce == _way1_hit_T_1 ? cache_data_206 : _GEN_1229; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1231 = 10'hcf == _way1_hit_T_1 ? cache_data_207 : _GEN_1230; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1232 = 10'hd0 == _way1_hit_T_1 ? cache_data_208 : _GEN_1231; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1233 = 10'hd1 == _way1_hit_T_1 ? cache_data_209 : _GEN_1232; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1234 = 10'hd2 == _way1_hit_T_1 ? cache_data_210 : _GEN_1233; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1235 = 10'hd3 == _way1_hit_T_1 ? cache_data_211 : _GEN_1234; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1236 = 10'hd4 == _way1_hit_T_1 ? cache_data_212 : _GEN_1235; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1237 = 10'hd5 == _way1_hit_T_1 ? cache_data_213 : _GEN_1236; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1238 = 10'hd6 == _way1_hit_T_1 ? cache_data_214 : _GEN_1237; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1239 = 10'hd7 == _way1_hit_T_1 ? cache_data_215 : _GEN_1238; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1240 = 10'hd8 == _way1_hit_T_1 ? cache_data_216 : _GEN_1239; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1241 = 10'hd9 == _way1_hit_T_1 ? cache_data_217 : _GEN_1240; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1242 = 10'hda == _way1_hit_T_1 ? cache_data_218 : _GEN_1241; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1243 = 10'hdb == _way1_hit_T_1 ? cache_data_219 : _GEN_1242; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1244 = 10'hdc == _way1_hit_T_1 ? cache_data_220 : _GEN_1243; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1245 = 10'hdd == _way1_hit_T_1 ? cache_data_221 : _GEN_1244; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1246 = 10'hde == _way1_hit_T_1 ? cache_data_222 : _GEN_1245; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1247 = 10'hdf == _way1_hit_T_1 ? cache_data_223 : _GEN_1246; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1248 = 10'he0 == _way1_hit_T_1 ? cache_data_224 : _GEN_1247; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1249 = 10'he1 == _way1_hit_T_1 ? cache_data_225 : _GEN_1248; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1250 = 10'he2 == _way1_hit_T_1 ? cache_data_226 : _GEN_1249; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1251 = 10'he3 == _way1_hit_T_1 ? cache_data_227 : _GEN_1250; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1252 = 10'he4 == _way1_hit_T_1 ? cache_data_228 : _GEN_1251; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1253 = 10'he5 == _way1_hit_T_1 ? cache_data_229 : _GEN_1252; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1254 = 10'he6 == _way1_hit_T_1 ? cache_data_230 : _GEN_1253; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1255 = 10'he7 == _way1_hit_T_1 ? cache_data_231 : _GEN_1254; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1256 = 10'he8 == _way1_hit_T_1 ? cache_data_232 : _GEN_1255; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1257 = 10'he9 == _way1_hit_T_1 ? cache_data_233 : _GEN_1256; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1258 = 10'hea == _way1_hit_T_1 ? cache_data_234 : _GEN_1257; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1259 = 10'heb == _way1_hit_T_1 ? cache_data_235 : _GEN_1258; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1260 = 10'hec == _way1_hit_T_1 ? cache_data_236 : _GEN_1259; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1261 = 10'hed == _way1_hit_T_1 ? cache_data_237 : _GEN_1260; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1262 = 10'hee == _way1_hit_T_1 ? cache_data_238 : _GEN_1261; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1263 = 10'hef == _way1_hit_T_1 ? cache_data_239 : _GEN_1262; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1264 = 10'hf0 == _way1_hit_T_1 ? cache_data_240 : _GEN_1263; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1265 = 10'hf1 == _way1_hit_T_1 ? cache_data_241 : _GEN_1264; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1266 = 10'hf2 == _way1_hit_T_1 ? cache_data_242 : _GEN_1265; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1267 = 10'hf3 == _way1_hit_T_1 ? cache_data_243 : _GEN_1266; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1268 = 10'hf4 == _way1_hit_T_1 ? cache_data_244 : _GEN_1267; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1269 = 10'hf5 == _way1_hit_T_1 ? cache_data_245 : _GEN_1268; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1270 = 10'hf6 == _way1_hit_T_1 ? cache_data_246 : _GEN_1269; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1271 = 10'hf7 == _way1_hit_T_1 ? cache_data_247 : _GEN_1270; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1272 = 10'hf8 == _way1_hit_T_1 ? cache_data_248 : _GEN_1271; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1273 = 10'hf9 == _way1_hit_T_1 ? cache_data_249 : _GEN_1272; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1274 = 10'hfa == _way1_hit_T_1 ? cache_data_250 : _GEN_1273; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1275 = 10'hfb == _way1_hit_T_1 ? cache_data_251 : _GEN_1274; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1276 = 10'hfc == _way1_hit_T_1 ? cache_data_252 : _GEN_1275; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1277 = 10'hfd == _way1_hit_T_1 ? cache_data_253 : _GEN_1276; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1278 = 10'hfe == _way1_hit_T_1 ? cache_data_254 : _GEN_1277; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1279 = 10'hff == _way1_hit_T_1 ? cache_data_255 : _GEN_1278; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1280 = 10'h100 == _way1_hit_T_1 ? cache_data_256 : _GEN_1279; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1281 = 10'h101 == _way1_hit_T_1 ? cache_data_257 : _GEN_1280; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1282 = 10'h102 == _way1_hit_T_1 ? cache_data_258 : _GEN_1281; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1283 = 10'h103 == _way1_hit_T_1 ? cache_data_259 : _GEN_1282; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1284 = 10'h104 == _way1_hit_T_1 ? cache_data_260 : _GEN_1283; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1285 = 10'h105 == _way1_hit_T_1 ? cache_data_261 : _GEN_1284; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1286 = 10'h106 == _way1_hit_T_1 ? cache_data_262 : _GEN_1285; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1287 = 10'h107 == _way1_hit_T_1 ? cache_data_263 : _GEN_1286; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1288 = 10'h108 == _way1_hit_T_1 ? cache_data_264 : _GEN_1287; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1289 = 10'h109 == _way1_hit_T_1 ? cache_data_265 : _GEN_1288; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1290 = 10'h10a == _way1_hit_T_1 ? cache_data_266 : _GEN_1289; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1291 = 10'h10b == _way1_hit_T_1 ? cache_data_267 : _GEN_1290; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1292 = 10'h10c == _way1_hit_T_1 ? cache_data_268 : _GEN_1291; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1293 = 10'h10d == _way1_hit_T_1 ? cache_data_269 : _GEN_1292; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1294 = 10'h10e == _way1_hit_T_1 ? cache_data_270 : _GEN_1293; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1295 = 10'h10f == _way1_hit_T_1 ? cache_data_271 : _GEN_1294; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1296 = 10'h110 == _way1_hit_T_1 ? cache_data_272 : _GEN_1295; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1297 = 10'h111 == _way1_hit_T_1 ? cache_data_273 : _GEN_1296; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1298 = 10'h112 == _way1_hit_T_1 ? cache_data_274 : _GEN_1297; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1299 = 10'h113 == _way1_hit_T_1 ? cache_data_275 : _GEN_1298; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1300 = 10'h114 == _way1_hit_T_1 ? cache_data_276 : _GEN_1299; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1301 = 10'h115 == _way1_hit_T_1 ? cache_data_277 : _GEN_1300; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1302 = 10'h116 == _way1_hit_T_1 ? cache_data_278 : _GEN_1301; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1303 = 10'h117 == _way1_hit_T_1 ? cache_data_279 : _GEN_1302; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1304 = 10'h118 == _way1_hit_T_1 ? cache_data_280 : _GEN_1303; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1305 = 10'h119 == _way1_hit_T_1 ? cache_data_281 : _GEN_1304; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1306 = 10'h11a == _way1_hit_T_1 ? cache_data_282 : _GEN_1305; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1307 = 10'h11b == _way1_hit_T_1 ? cache_data_283 : _GEN_1306; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1308 = 10'h11c == _way1_hit_T_1 ? cache_data_284 : _GEN_1307; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1309 = 10'h11d == _way1_hit_T_1 ? cache_data_285 : _GEN_1308; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1310 = 10'h11e == _way1_hit_T_1 ? cache_data_286 : _GEN_1309; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1311 = 10'h11f == _way1_hit_T_1 ? cache_data_287 : _GEN_1310; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1312 = 10'h120 == _way1_hit_T_1 ? cache_data_288 : _GEN_1311; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1313 = 10'h121 == _way1_hit_T_1 ? cache_data_289 : _GEN_1312; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1314 = 10'h122 == _way1_hit_T_1 ? cache_data_290 : _GEN_1313; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1315 = 10'h123 == _way1_hit_T_1 ? cache_data_291 : _GEN_1314; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1316 = 10'h124 == _way1_hit_T_1 ? cache_data_292 : _GEN_1315; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1317 = 10'h125 == _way1_hit_T_1 ? cache_data_293 : _GEN_1316; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1318 = 10'h126 == _way1_hit_T_1 ? cache_data_294 : _GEN_1317; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1319 = 10'h127 == _way1_hit_T_1 ? cache_data_295 : _GEN_1318; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1320 = 10'h128 == _way1_hit_T_1 ? cache_data_296 : _GEN_1319; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1321 = 10'h129 == _way1_hit_T_1 ? cache_data_297 : _GEN_1320; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1322 = 10'h12a == _way1_hit_T_1 ? cache_data_298 : _GEN_1321; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1323 = 10'h12b == _way1_hit_T_1 ? cache_data_299 : _GEN_1322; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1324 = 10'h12c == _way1_hit_T_1 ? cache_data_300 : _GEN_1323; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1325 = 10'h12d == _way1_hit_T_1 ? cache_data_301 : _GEN_1324; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1326 = 10'h12e == _way1_hit_T_1 ? cache_data_302 : _GEN_1325; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1327 = 10'h12f == _way1_hit_T_1 ? cache_data_303 : _GEN_1326; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1328 = 10'h130 == _way1_hit_T_1 ? cache_data_304 : _GEN_1327; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1329 = 10'h131 == _way1_hit_T_1 ? cache_data_305 : _GEN_1328; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1330 = 10'h132 == _way1_hit_T_1 ? cache_data_306 : _GEN_1329; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1331 = 10'h133 == _way1_hit_T_1 ? cache_data_307 : _GEN_1330; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1332 = 10'h134 == _way1_hit_T_1 ? cache_data_308 : _GEN_1331; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1333 = 10'h135 == _way1_hit_T_1 ? cache_data_309 : _GEN_1332; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1334 = 10'h136 == _way1_hit_T_1 ? cache_data_310 : _GEN_1333; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1335 = 10'h137 == _way1_hit_T_1 ? cache_data_311 : _GEN_1334; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1336 = 10'h138 == _way1_hit_T_1 ? cache_data_312 : _GEN_1335; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1337 = 10'h139 == _way1_hit_T_1 ? cache_data_313 : _GEN_1336; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1338 = 10'h13a == _way1_hit_T_1 ? cache_data_314 : _GEN_1337; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1339 = 10'h13b == _way1_hit_T_1 ? cache_data_315 : _GEN_1338; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1340 = 10'h13c == _way1_hit_T_1 ? cache_data_316 : _GEN_1339; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1341 = 10'h13d == _way1_hit_T_1 ? cache_data_317 : _GEN_1340; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1342 = 10'h13e == _way1_hit_T_1 ? cache_data_318 : _GEN_1341; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1343 = 10'h13f == _way1_hit_T_1 ? cache_data_319 : _GEN_1342; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1344 = 10'h140 == _way1_hit_T_1 ? cache_data_320 : _GEN_1343; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1345 = 10'h141 == _way1_hit_T_1 ? cache_data_321 : _GEN_1344; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1346 = 10'h142 == _way1_hit_T_1 ? cache_data_322 : _GEN_1345; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1347 = 10'h143 == _way1_hit_T_1 ? cache_data_323 : _GEN_1346; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1348 = 10'h144 == _way1_hit_T_1 ? cache_data_324 : _GEN_1347; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1349 = 10'h145 == _way1_hit_T_1 ? cache_data_325 : _GEN_1348; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1350 = 10'h146 == _way1_hit_T_1 ? cache_data_326 : _GEN_1349; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1351 = 10'h147 == _way1_hit_T_1 ? cache_data_327 : _GEN_1350; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1352 = 10'h148 == _way1_hit_T_1 ? cache_data_328 : _GEN_1351; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1353 = 10'h149 == _way1_hit_T_1 ? cache_data_329 : _GEN_1352; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1354 = 10'h14a == _way1_hit_T_1 ? cache_data_330 : _GEN_1353; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1355 = 10'h14b == _way1_hit_T_1 ? cache_data_331 : _GEN_1354; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1356 = 10'h14c == _way1_hit_T_1 ? cache_data_332 : _GEN_1355; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1357 = 10'h14d == _way1_hit_T_1 ? cache_data_333 : _GEN_1356; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1358 = 10'h14e == _way1_hit_T_1 ? cache_data_334 : _GEN_1357; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1359 = 10'h14f == _way1_hit_T_1 ? cache_data_335 : _GEN_1358; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1360 = 10'h150 == _way1_hit_T_1 ? cache_data_336 : _GEN_1359; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1361 = 10'h151 == _way1_hit_T_1 ? cache_data_337 : _GEN_1360; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1362 = 10'h152 == _way1_hit_T_1 ? cache_data_338 : _GEN_1361; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1363 = 10'h153 == _way1_hit_T_1 ? cache_data_339 : _GEN_1362; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1364 = 10'h154 == _way1_hit_T_1 ? cache_data_340 : _GEN_1363; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1365 = 10'h155 == _way1_hit_T_1 ? cache_data_341 : _GEN_1364; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1366 = 10'h156 == _way1_hit_T_1 ? cache_data_342 : _GEN_1365; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1367 = 10'h157 == _way1_hit_T_1 ? cache_data_343 : _GEN_1366; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1368 = 10'h158 == _way1_hit_T_1 ? cache_data_344 : _GEN_1367; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1369 = 10'h159 == _way1_hit_T_1 ? cache_data_345 : _GEN_1368; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1370 = 10'h15a == _way1_hit_T_1 ? cache_data_346 : _GEN_1369; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1371 = 10'h15b == _way1_hit_T_1 ? cache_data_347 : _GEN_1370; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1372 = 10'h15c == _way1_hit_T_1 ? cache_data_348 : _GEN_1371; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1373 = 10'h15d == _way1_hit_T_1 ? cache_data_349 : _GEN_1372; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1374 = 10'h15e == _way1_hit_T_1 ? cache_data_350 : _GEN_1373; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1375 = 10'h15f == _way1_hit_T_1 ? cache_data_351 : _GEN_1374; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1376 = 10'h160 == _way1_hit_T_1 ? cache_data_352 : _GEN_1375; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1377 = 10'h161 == _way1_hit_T_1 ? cache_data_353 : _GEN_1376; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1378 = 10'h162 == _way1_hit_T_1 ? cache_data_354 : _GEN_1377; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1379 = 10'h163 == _way1_hit_T_1 ? cache_data_355 : _GEN_1378; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1380 = 10'h164 == _way1_hit_T_1 ? cache_data_356 : _GEN_1379; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1381 = 10'h165 == _way1_hit_T_1 ? cache_data_357 : _GEN_1380; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1382 = 10'h166 == _way1_hit_T_1 ? cache_data_358 : _GEN_1381; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1383 = 10'h167 == _way1_hit_T_1 ? cache_data_359 : _GEN_1382; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1384 = 10'h168 == _way1_hit_T_1 ? cache_data_360 : _GEN_1383; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1385 = 10'h169 == _way1_hit_T_1 ? cache_data_361 : _GEN_1384; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1386 = 10'h16a == _way1_hit_T_1 ? cache_data_362 : _GEN_1385; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1387 = 10'h16b == _way1_hit_T_1 ? cache_data_363 : _GEN_1386; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1388 = 10'h16c == _way1_hit_T_1 ? cache_data_364 : _GEN_1387; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1389 = 10'h16d == _way1_hit_T_1 ? cache_data_365 : _GEN_1388; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1390 = 10'h16e == _way1_hit_T_1 ? cache_data_366 : _GEN_1389; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1391 = 10'h16f == _way1_hit_T_1 ? cache_data_367 : _GEN_1390; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1392 = 10'h170 == _way1_hit_T_1 ? cache_data_368 : _GEN_1391; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1393 = 10'h171 == _way1_hit_T_1 ? cache_data_369 : _GEN_1392; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1394 = 10'h172 == _way1_hit_T_1 ? cache_data_370 : _GEN_1393; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1395 = 10'h173 == _way1_hit_T_1 ? cache_data_371 : _GEN_1394; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1396 = 10'h174 == _way1_hit_T_1 ? cache_data_372 : _GEN_1395; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1397 = 10'h175 == _way1_hit_T_1 ? cache_data_373 : _GEN_1396; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1398 = 10'h176 == _way1_hit_T_1 ? cache_data_374 : _GEN_1397; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1399 = 10'h177 == _way1_hit_T_1 ? cache_data_375 : _GEN_1398; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1400 = 10'h178 == _way1_hit_T_1 ? cache_data_376 : _GEN_1399; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1401 = 10'h179 == _way1_hit_T_1 ? cache_data_377 : _GEN_1400; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1402 = 10'h17a == _way1_hit_T_1 ? cache_data_378 : _GEN_1401; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1403 = 10'h17b == _way1_hit_T_1 ? cache_data_379 : _GEN_1402; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1404 = 10'h17c == _way1_hit_T_1 ? cache_data_380 : _GEN_1403; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1405 = 10'h17d == _way1_hit_T_1 ? cache_data_381 : _GEN_1404; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1406 = 10'h17e == _way1_hit_T_1 ? cache_data_382 : _GEN_1405; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1407 = 10'h17f == _way1_hit_T_1 ? cache_data_383 : _GEN_1406; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1408 = 10'h180 == _way1_hit_T_1 ? cache_data_384 : _GEN_1407; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1409 = 10'h181 == _way1_hit_T_1 ? cache_data_385 : _GEN_1408; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1410 = 10'h182 == _way1_hit_T_1 ? cache_data_386 : _GEN_1409; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1411 = 10'h183 == _way1_hit_T_1 ? cache_data_387 : _GEN_1410; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1412 = 10'h184 == _way1_hit_T_1 ? cache_data_388 : _GEN_1411; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1413 = 10'h185 == _way1_hit_T_1 ? cache_data_389 : _GEN_1412; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1414 = 10'h186 == _way1_hit_T_1 ? cache_data_390 : _GEN_1413; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1415 = 10'h187 == _way1_hit_T_1 ? cache_data_391 : _GEN_1414; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1416 = 10'h188 == _way1_hit_T_1 ? cache_data_392 : _GEN_1415; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1417 = 10'h189 == _way1_hit_T_1 ? cache_data_393 : _GEN_1416; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1418 = 10'h18a == _way1_hit_T_1 ? cache_data_394 : _GEN_1417; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1419 = 10'h18b == _way1_hit_T_1 ? cache_data_395 : _GEN_1418; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1420 = 10'h18c == _way1_hit_T_1 ? cache_data_396 : _GEN_1419; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1421 = 10'h18d == _way1_hit_T_1 ? cache_data_397 : _GEN_1420; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1422 = 10'h18e == _way1_hit_T_1 ? cache_data_398 : _GEN_1421; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1423 = 10'h18f == _way1_hit_T_1 ? cache_data_399 : _GEN_1422; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1424 = 10'h190 == _way1_hit_T_1 ? cache_data_400 : _GEN_1423; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1425 = 10'h191 == _way1_hit_T_1 ? cache_data_401 : _GEN_1424; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1426 = 10'h192 == _way1_hit_T_1 ? cache_data_402 : _GEN_1425; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1427 = 10'h193 == _way1_hit_T_1 ? cache_data_403 : _GEN_1426; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1428 = 10'h194 == _way1_hit_T_1 ? cache_data_404 : _GEN_1427; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1429 = 10'h195 == _way1_hit_T_1 ? cache_data_405 : _GEN_1428; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1430 = 10'h196 == _way1_hit_T_1 ? cache_data_406 : _GEN_1429; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1431 = 10'h197 == _way1_hit_T_1 ? cache_data_407 : _GEN_1430; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1432 = 10'h198 == _way1_hit_T_1 ? cache_data_408 : _GEN_1431; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1433 = 10'h199 == _way1_hit_T_1 ? cache_data_409 : _GEN_1432; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1434 = 10'h19a == _way1_hit_T_1 ? cache_data_410 : _GEN_1433; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1435 = 10'h19b == _way1_hit_T_1 ? cache_data_411 : _GEN_1434; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1436 = 10'h19c == _way1_hit_T_1 ? cache_data_412 : _GEN_1435; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1437 = 10'h19d == _way1_hit_T_1 ? cache_data_413 : _GEN_1436; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1438 = 10'h19e == _way1_hit_T_1 ? cache_data_414 : _GEN_1437; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1439 = 10'h19f == _way1_hit_T_1 ? cache_data_415 : _GEN_1438; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1440 = 10'h1a0 == _way1_hit_T_1 ? cache_data_416 : _GEN_1439; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1441 = 10'h1a1 == _way1_hit_T_1 ? cache_data_417 : _GEN_1440; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1442 = 10'h1a2 == _way1_hit_T_1 ? cache_data_418 : _GEN_1441; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1443 = 10'h1a3 == _way1_hit_T_1 ? cache_data_419 : _GEN_1442; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1444 = 10'h1a4 == _way1_hit_T_1 ? cache_data_420 : _GEN_1443; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1445 = 10'h1a5 == _way1_hit_T_1 ? cache_data_421 : _GEN_1444; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1446 = 10'h1a6 == _way1_hit_T_1 ? cache_data_422 : _GEN_1445; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1447 = 10'h1a7 == _way1_hit_T_1 ? cache_data_423 : _GEN_1446; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1448 = 10'h1a8 == _way1_hit_T_1 ? cache_data_424 : _GEN_1447; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1449 = 10'h1a9 == _way1_hit_T_1 ? cache_data_425 : _GEN_1448; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1450 = 10'h1aa == _way1_hit_T_1 ? cache_data_426 : _GEN_1449; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1451 = 10'h1ab == _way1_hit_T_1 ? cache_data_427 : _GEN_1450; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1452 = 10'h1ac == _way1_hit_T_1 ? cache_data_428 : _GEN_1451; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1453 = 10'h1ad == _way1_hit_T_1 ? cache_data_429 : _GEN_1452; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1454 = 10'h1ae == _way1_hit_T_1 ? cache_data_430 : _GEN_1453; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1455 = 10'h1af == _way1_hit_T_1 ? cache_data_431 : _GEN_1454; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1456 = 10'h1b0 == _way1_hit_T_1 ? cache_data_432 : _GEN_1455; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1457 = 10'h1b1 == _way1_hit_T_1 ? cache_data_433 : _GEN_1456; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1458 = 10'h1b2 == _way1_hit_T_1 ? cache_data_434 : _GEN_1457; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1459 = 10'h1b3 == _way1_hit_T_1 ? cache_data_435 : _GEN_1458; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1460 = 10'h1b4 == _way1_hit_T_1 ? cache_data_436 : _GEN_1459; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1461 = 10'h1b5 == _way1_hit_T_1 ? cache_data_437 : _GEN_1460; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1462 = 10'h1b6 == _way1_hit_T_1 ? cache_data_438 : _GEN_1461; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1463 = 10'h1b7 == _way1_hit_T_1 ? cache_data_439 : _GEN_1462; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1464 = 10'h1b8 == _way1_hit_T_1 ? cache_data_440 : _GEN_1463; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1465 = 10'h1b9 == _way1_hit_T_1 ? cache_data_441 : _GEN_1464; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1466 = 10'h1ba == _way1_hit_T_1 ? cache_data_442 : _GEN_1465; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1467 = 10'h1bb == _way1_hit_T_1 ? cache_data_443 : _GEN_1466; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1468 = 10'h1bc == _way1_hit_T_1 ? cache_data_444 : _GEN_1467; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1469 = 10'h1bd == _way1_hit_T_1 ? cache_data_445 : _GEN_1468; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1470 = 10'h1be == _way1_hit_T_1 ? cache_data_446 : _GEN_1469; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1471 = 10'h1bf == _way1_hit_T_1 ? cache_data_447 : _GEN_1470; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1472 = 10'h1c0 == _way1_hit_T_1 ? cache_data_448 : _GEN_1471; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1473 = 10'h1c1 == _way1_hit_T_1 ? cache_data_449 : _GEN_1472; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1474 = 10'h1c2 == _way1_hit_T_1 ? cache_data_450 : _GEN_1473; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1475 = 10'h1c3 == _way1_hit_T_1 ? cache_data_451 : _GEN_1474; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1476 = 10'h1c4 == _way1_hit_T_1 ? cache_data_452 : _GEN_1475; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1477 = 10'h1c5 == _way1_hit_T_1 ? cache_data_453 : _GEN_1476; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1478 = 10'h1c6 == _way1_hit_T_1 ? cache_data_454 : _GEN_1477; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1479 = 10'h1c7 == _way1_hit_T_1 ? cache_data_455 : _GEN_1478; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1480 = 10'h1c8 == _way1_hit_T_1 ? cache_data_456 : _GEN_1479; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1481 = 10'h1c9 == _way1_hit_T_1 ? cache_data_457 : _GEN_1480; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1482 = 10'h1ca == _way1_hit_T_1 ? cache_data_458 : _GEN_1481; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1483 = 10'h1cb == _way1_hit_T_1 ? cache_data_459 : _GEN_1482; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1484 = 10'h1cc == _way1_hit_T_1 ? cache_data_460 : _GEN_1483; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1485 = 10'h1cd == _way1_hit_T_1 ? cache_data_461 : _GEN_1484; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1486 = 10'h1ce == _way1_hit_T_1 ? cache_data_462 : _GEN_1485; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1487 = 10'h1cf == _way1_hit_T_1 ? cache_data_463 : _GEN_1486; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1488 = 10'h1d0 == _way1_hit_T_1 ? cache_data_464 : _GEN_1487; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1489 = 10'h1d1 == _way1_hit_T_1 ? cache_data_465 : _GEN_1488; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1490 = 10'h1d2 == _way1_hit_T_1 ? cache_data_466 : _GEN_1489; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1491 = 10'h1d3 == _way1_hit_T_1 ? cache_data_467 : _GEN_1490; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1492 = 10'h1d4 == _way1_hit_T_1 ? cache_data_468 : _GEN_1491; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1493 = 10'h1d5 == _way1_hit_T_1 ? cache_data_469 : _GEN_1492; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1494 = 10'h1d6 == _way1_hit_T_1 ? cache_data_470 : _GEN_1493; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1495 = 10'h1d7 == _way1_hit_T_1 ? cache_data_471 : _GEN_1494; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1496 = 10'h1d8 == _way1_hit_T_1 ? cache_data_472 : _GEN_1495; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1497 = 10'h1d9 == _way1_hit_T_1 ? cache_data_473 : _GEN_1496; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1498 = 10'h1da == _way1_hit_T_1 ? cache_data_474 : _GEN_1497; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1499 = 10'h1db == _way1_hit_T_1 ? cache_data_475 : _GEN_1498; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1500 = 10'h1dc == _way1_hit_T_1 ? cache_data_476 : _GEN_1499; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1501 = 10'h1dd == _way1_hit_T_1 ? cache_data_477 : _GEN_1500; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1502 = 10'h1de == _way1_hit_T_1 ? cache_data_478 : _GEN_1501; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1503 = 10'h1df == _way1_hit_T_1 ? cache_data_479 : _GEN_1502; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1504 = 10'h1e0 == _way1_hit_T_1 ? cache_data_480 : _GEN_1503; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1505 = 10'h1e1 == _way1_hit_T_1 ? cache_data_481 : _GEN_1504; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1506 = 10'h1e2 == _way1_hit_T_1 ? cache_data_482 : _GEN_1505; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1507 = 10'h1e3 == _way1_hit_T_1 ? cache_data_483 : _GEN_1506; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1508 = 10'h1e4 == _way1_hit_T_1 ? cache_data_484 : _GEN_1507; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1509 = 10'h1e5 == _way1_hit_T_1 ? cache_data_485 : _GEN_1508; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1510 = 10'h1e6 == _way1_hit_T_1 ? cache_data_486 : _GEN_1509; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1511 = 10'h1e7 == _way1_hit_T_1 ? cache_data_487 : _GEN_1510; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1512 = 10'h1e8 == _way1_hit_T_1 ? cache_data_488 : _GEN_1511; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1513 = 10'h1e9 == _way1_hit_T_1 ? cache_data_489 : _GEN_1512; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1514 = 10'h1ea == _way1_hit_T_1 ? cache_data_490 : _GEN_1513; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1515 = 10'h1eb == _way1_hit_T_1 ? cache_data_491 : _GEN_1514; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1516 = 10'h1ec == _way1_hit_T_1 ? cache_data_492 : _GEN_1515; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1517 = 10'h1ed == _way1_hit_T_1 ? cache_data_493 : _GEN_1516; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1518 = 10'h1ee == _way1_hit_T_1 ? cache_data_494 : _GEN_1517; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1519 = 10'h1ef == _way1_hit_T_1 ? cache_data_495 : _GEN_1518; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1520 = 10'h1f0 == _way1_hit_T_1 ? cache_data_496 : _GEN_1519; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1521 = 10'h1f1 == _way1_hit_T_1 ? cache_data_497 : _GEN_1520; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1522 = 10'h1f2 == _way1_hit_T_1 ? cache_data_498 : _GEN_1521; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1523 = 10'h1f3 == _way1_hit_T_1 ? cache_data_499 : _GEN_1522; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1524 = 10'h1f4 == _way1_hit_T_1 ? cache_data_500 : _GEN_1523; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1525 = 10'h1f5 == _way1_hit_T_1 ? cache_data_501 : _GEN_1524; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1526 = 10'h1f6 == _way1_hit_T_1 ? cache_data_502 : _GEN_1525; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1527 = 10'h1f7 == _way1_hit_T_1 ? cache_data_503 : _GEN_1526; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1528 = 10'h1f8 == _way1_hit_T_1 ? cache_data_504 : _GEN_1527; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1529 = 10'h1f9 == _way1_hit_T_1 ? cache_data_505 : _GEN_1528; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1530 = 10'h1fa == _way1_hit_T_1 ? cache_data_506 : _GEN_1529; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1531 = 10'h1fb == _way1_hit_T_1 ? cache_data_507 : _GEN_1530; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1532 = 10'h1fc == _way1_hit_T_1 ? cache_data_508 : _GEN_1531; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1533 = 10'h1fd == _way1_hit_T_1 ? cache_data_509 : _GEN_1532; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1534 = 10'h1fe == _way1_hit_T_1 ? cache_data_510 : _GEN_1533; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1535 = 10'h1ff == _way1_hit_T_1 ? cache_data_511 : _GEN_1534; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1536 = 10'h200 == _way1_hit_T_1 ? cache_data_512 : _GEN_1535; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1537 = 10'h201 == _way1_hit_T_1 ? cache_data_513 : _GEN_1536; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1538 = 10'h202 == _way1_hit_T_1 ? cache_data_514 : _GEN_1537; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1539 = 10'h203 == _way1_hit_T_1 ? cache_data_515 : _GEN_1538; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1540 = 10'h204 == _way1_hit_T_1 ? cache_data_516 : _GEN_1539; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1541 = 10'h205 == _way1_hit_T_1 ? cache_data_517 : _GEN_1540; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1542 = 10'h206 == _way1_hit_T_1 ? cache_data_518 : _GEN_1541; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1543 = 10'h207 == _way1_hit_T_1 ? cache_data_519 : _GEN_1542; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1544 = 10'h208 == _way1_hit_T_1 ? cache_data_520 : _GEN_1543; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1545 = 10'h209 == _way1_hit_T_1 ? cache_data_521 : _GEN_1544; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1546 = 10'h20a == _way1_hit_T_1 ? cache_data_522 : _GEN_1545; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1547 = 10'h20b == _way1_hit_T_1 ? cache_data_523 : _GEN_1546; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1548 = 10'h20c == _way1_hit_T_1 ? cache_data_524 : _GEN_1547; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1549 = 10'h20d == _way1_hit_T_1 ? cache_data_525 : _GEN_1548; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1550 = 10'h20e == _way1_hit_T_1 ? cache_data_526 : _GEN_1549; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1551 = 10'h20f == _way1_hit_T_1 ? cache_data_527 : _GEN_1550; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1552 = 10'h210 == _way1_hit_T_1 ? cache_data_528 : _GEN_1551; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1553 = 10'h211 == _way1_hit_T_1 ? cache_data_529 : _GEN_1552; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1554 = 10'h212 == _way1_hit_T_1 ? cache_data_530 : _GEN_1553; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1555 = 10'h213 == _way1_hit_T_1 ? cache_data_531 : _GEN_1554; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1556 = 10'h214 == _way1_hit_T_1 ? cache_data_532 : _GEN_1555; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1557 = 10'h215 == _way1_hit_T_1 ? cache_data_533 : _GEN_1556; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1558 = 10'h216 == _way1_hit_T_1 ? cache_data_534 : _GEN_1557; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1559 = 10'h217 == _way1_hit_T_1 ? cache_data_535 : _GEN_1558; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1560 = 10'h218 == _way1_hit_T_1 ? cache_data_536 : _GEN_1559; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1561 = 10'h219 == _way1_hit_T_1 ? cache_data_537 : _GEN_1560; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1562 = 10'h21a == _way1_hit_T_1 ? cache_data_538 : _GEN_1561; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1563 = 10'h21b == _way1_hit_T_1 ? cache_data_539 : _GEN_1562; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1564 = 10'h21c == _way1_hit_T_1 ? cache_data_540 : _GEN_1563; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1565 = 10'h21d == _way1_hit_T_1 ? cache_data_541 : _GEN_1564; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1566 = 10'h21e == _way1_hit_T_1 ? cache_data_542 : _GEN_1565; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1567 = 10'h21f == _way1_hit_T_1 ? cache_data_543 : _GEN_1566; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1568 = 10'h220 == _way1_hit_T_1 ? cache_data_544 : _GEN_1567; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1569 = 10'h221 == _way1_hit_T_1 ? cache_data_545 : _GEN_1568; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1570 = 10'h222 == _way1_hit_T_1 ? cache_data_546 : _GEN_1569; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1571 = 10'h223 == _way1_hit_T_1 ? cache_data_547 : _GEN_1570; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1572 = 10'h224 == _way1_hit_T_1 ? cache_data_548 : _GEN_1571; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1573 = 10'h225 == _way1_hit_T_1 ? cache_data_549 : _GEN_1572; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1574 = 10'h226 == _way1_hit_T_1 ? cache_data_550 : _GEN_1573; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1575 = 10'h227 == _way1_hit_T_1 ? cache_data_551 : _GEN_1574; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1576 = 10'h228 == _way1_hit_T_1 ? cache_data_552 : _GEN_1575; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1577 = 10'h229 == _way1_hit_T_1 ? cache_data_553 : _GEN_1576; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1578 = 10'h22a == _way1_hit_T_1 ? cache_data_554 : _GEN_1577; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1579 = 10'h22b == _way1_hit_T_1 ? cache_data_555 : _GEN_1578; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1580 = 10'h22c == _way1_hit_T_1 ? cache_data_556 : _GEN_1579; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1581 = 10'h22d == _way1_hit_T_1 ? cache_data_557 : _GEN_1580; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1582 = 10'h22e == _way1_hit_T_1 ? cache_data_558 : _GEN_1581; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1583 = 10'h22f == _way1_hit_T_1 ? cache_data_559 : _GEN_1582; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1584 = 10'h230 == _way1_hit_T_1 ? cache_data_560 : _GEN_1583; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1585 = 10'h231 == _way1_hit_T_1 ? cache_data_561 : _GEN_1584; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1586 = 10'h232 == _way1_hit_T_1 ? cache_data_562 : _GEN_1585; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1587 = 10'h233 == _way1_hit_T_1 ? cache_data_563 : _GEN_1586; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1588 = 10'h234 == _way1_hit_T_1 ? cache_data_564 : _GEN_1587; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1589 = 10'h235 == _way1_hit_T_1 ? cache_data_565 : _GEN_1588; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1590 = 10'h236 == _way1_hit_T_1 ? cache_data_566 : _GEN_1589; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1591 = 10'h237 == _way1_hit_T_1 ? cache_data_567 : _GEN_1590; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1592 = 10'h238 == _way1_hit_T_1 ? cache_data_568 : _GEN_1591; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1593 = 10'h239 == _way1_hit_T_1 ? cache_data_569 : _GEN_1592; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1594 = 10'h23a == _way1_hit_T_1 ? cache_data_570 : _GEN_1593; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1595 = 10'h23b == _way1_hit_T_1 ? cache_data_571 : _GEN_1594; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1596 = 10'h23c == _way1_hit_T_1 ? cache_data_572 : _GEN_1595; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1597 = 10'h23d == _way1_hit_T_1 ? cache_data_573 : _GEN_1596; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1598 = 10'h23e == _way1_hit_T_1 ? cache_data_574 : _GEN_1597; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1599 = 10'h23f == _way1_hit_T_1 ? cache_data_575 : _GEN_1598; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1600 = 10'h240 == _way1_hit_T_1 ? cache_data_576 : _GEN_1599; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1601 = 10'h241 == _way1_hit_T_1 ? cache_data_577 : _GEN_1600; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1602 = 10'h242 == _way1_hit_T_1 ? cache_data_578 : _GEN_1601; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1603 = 10'h243 == _way1_hit_T_1 ? cache_data_579 : _GEN_1602; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1604 = 10'h244 == _way1_hit_T_1 ? cache_data_580 : _GEN_1603; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1605 = 10'h245 == _way1_hit_T_1 ? cache_data_581 : _GEN_1604; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1606 = 10'h246 == _way1_hit_T_1 ? cache_data_582 : _GEN_1605; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1607 = 10'h247 == _way1_hit_T_1 ? cache_data_583 : _GEN_1606; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1608 = 10'h248 == _way1_hit_T_1 ? cache_data_584 : _GEN_1607; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1609 = 10'h249 == _way1_hit_T_1 ? cache_data_585 : _GEN_1608; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1610 = 10'h24a == _way1_hit_T_1 ? cache_data_586 : _GEN_1609; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1611 = 10'h24b == _way1_hit_T_1 ? cache_data_587 : _GEN_1610; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1612 = 10'h24c == _way1_hit_T_1 ? cache_data_588 : _GEN_1611; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1613 = 10'h24d == _way1_hit_T_1 ? cache_data_589 : _GEN_1612; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1614 = 10'h24e == _way1_hit_T_1 ? cache_data_590 : _GEN_1613; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1615 = 10'h24f == _way1_hit_T_1 ? cache_data_591 : _GEN_1614; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1616 = 10'h250 == _way1_hit_T_1 ? cache_data_592 : _GEN_1615; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1617 = 10'h251 == _way1_hit_T_1 ? cache_data_593 : _GEN_1616; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1618 = 10'h252 == _way1_hit_T_1 ? cache_data_594 : _GEN_1617; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1619 = 10'h253 == _way1_hit_T_1 ? cache_data_595 : _GEN_1618; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1620 = 10'h254 == _way1_hit_T_1 ? cache_data_596 : _GEN_1619; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1621 = 10'h255 == _way1_hit_T_1 ? cache_data_597 : _GEN_1620; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1622 = 10'h256 == _way1_hit_T_1 ? cache_data_598 : _GEN_1621; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1623 = 10'h257 == _way1_hit_T_1 ? cache_data_599 : _GEN_1622; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1624 = 10'h258 == _way1_hit_T_1 ? cache_data_600 : _GEN_1623; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1625 = 10'h259 == _way1_hit_T_1 ? cache_data_601 : _GEN_1624; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1626 = 10'h25a == _way1_hit_T_1 ? cache_data_602 : _GEN_1625; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1627 = 10'h25b == _way1_hit_T_1 ? cache_data_603 : _GEN_1626; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1628 = 10'h25c == _way1_hit_T_1 ? cache_data_604 : _GEN_1627; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1629 = 10'h25d == _way1_hit_T_1 ? cache_data_605 : _GEN_1628; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1630 = 10'h25e == _way1_hit_T_1 ? cache_data_606 : _GEN_1629; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1631 = 10'h25f == _way1_hit_T_1 ? cache_data_607 : _GEN_1630; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1632 = 10'h260 == _way1_hit_T_1 ? cache_data_608 : _GEN_1631; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1633 = 10'h261 == _way1_hit_T_1 ? cache_data_609 : _GEN_1632; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1634 = 10'h262 == _way1_hit_T_1 ? cache_data_610 : _GEN_1633; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1635 = 10'h263 == _way1_hit_T_1 ? cache_data_611 : _GEN_1634; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1636 = 10'h264 == _way1_hit_T_1 ? cache_data_612 : _GEN_1635; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1637 = 10'h265 == _way1_hit_T_1 ? cache_data_613 : _GEN_1636; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1638 = 10'h266 == _way1_hit_T_1 ? cache_data_614 : _GEN_1637; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1639 = 10'h267 == _way1_hit_T_1 ? cache_data_615 : _GEN_1638; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1640 = 10'h268 == _way1_hit_T_1 ? cache_data_616 : _GEN_1639; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1641 = 10'h269 == _way1_hit_T_1 ? cache_data_617 : _GEN_1640; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1642 = 10'h26a == _way1_hit_T_1 ? cache_data_618 : _GEN_1641; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1643 = 10'h26b == _way1_hit_T_1 ? cache_data_619 : _GEN_1642; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1644 = 10'h26c == _way1_hit_T_1 ? cache_data_620 : _GEN_1643; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1645 = 10'h26d == _way1_hit_T_1 ? cache_data_621 : _GEN_1644; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1646 = 10'h26e == _way1_hit_T_1 ? cache_data_622 : _GEN_1645; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1647 = 10'h26f == _way1_hit_T_1 ? cache_data_623 : _GEN_1646; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1648 = 10'h270 == _way1_hit_T_1 ? cache_data_624 : _GEN_1647; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1649 = 10'h271 == _way1_hit_T_1 ? cache_data_625 : _GEN_1648; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1650 = 10'h272 == _way1_hit_T_1 ? cache_data_626 : _GEN_1649; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1651 = 10'h273 == _way1_hit_T_1 ? cache_data_627 : _GEN_1650; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1652 = 10'h274 == _way1_hit_T_1 ? cache_data_628 : _GEN_1651; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1653 = 10'h275 == _way1_hit_T_1 ? cache_data_629 : _GEN_1652; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1654 = 10'h276 == _way1_hit_T_1 ? cache_data_630 : _GEN_1653; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1655 = 10'h277 == _way1_hit_T_1 ? cache_data_631 : _GEN_1654; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1656 = 10'h278 == _way1_hit_T_1 ? cache_data_632 : _GEN_1655; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1657 = 10'h279 == _way1_hit_T_1 ? cache_data_633 : _GEN_1656; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1658 = 10'h27a == _way1_hit_T_1 ? cache_data_634 : _GEN_1657; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1659 = 10'h27b == _way1_hit_T_1 ? cache_data_635 : _GEN_1658; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1660 = 10'h27c == _way1_hit_T_1 ? cache_data_636 : _GEN_1659; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1661 = 10'h27d == _way1_hit_T_1 ? cache_data_637 : _GEN_1660; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1662 = 10'h27e == _way1_hit_T_1 ? cache_data_638 : _GEN_1661; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1663 = 10'h27f == _way1_hit_T_1 ? cache_data_639 : _GEN_1662; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1664 = 10'h280 == _way1_hit_T_1 ? cache_data_640 : _GEN_1663; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1665 = 10'h281 == _way1_hit_T_1 ? cache_data_641 : _GEN_1664; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1666 = 10'h282 == _way1_hit_T_1 ? cache_data_642 : _GEN_1665; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1667 = 10'h283 == _way1_hit_T_1 ? cache_data_643 : _GEN_1666; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1668 = 10'h284 == _way1_hit_T_1 ? cache_data_644 : _GEN_1667; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1669 = 10'h285 == _way1_hit_T_1 ? cache_data_645 : _GEN_1668; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1670 = 10'h286 == _way1_hit_T_1 ? cache_data_646 : _GEN_1669; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1671 = 10'h287 == _way1_hit_T_1 ? cache_data_647 : _GEN_1670; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1672 = 10'h288 == _way1_hit_T_1 ? cache_data_648 : _GEN_1671; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1673 = 10'h289 == _way1_hit_T_1 ? cache_data_649 : _GEN_1672; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1674 = 10'h28a == _way1_hit_T_1 ? cache_data_650 : _GEN_1673; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1675 = 10'h28b == _way1_hit_T_1 ? cache_data_651 : _GEN_1674; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1676 = 10'h28c == _way1_hit_T_1 ? cache_data_652 : _GEN_1675; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1677 = 10'h28d == _way1_hit_T_1 ? cache_data_653 : _GEN_1676; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1678 = 10'h28e == _way1_hit_T_1 ? cache_data_654 : _GEN_1677; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1679 = 10'h28f == _way1_hit_T_1 ? cache_data_655 : _GEN_1678; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1680 = 10'h290 == _way1_hit_T_1 ? cache_data_656 : _GEN_1679; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1681 = 10'h291 == _way1_hit_T_1 ? cache_data_657 : _GEN_1680; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1682 = 10'h292 == _way1_hit_T_1 ? cache_data_658 : _GEN_1681; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1683 = 10'h293 == _way1_hit_T_1 ? cache_data_659 : _GEN_1682; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1684 = 10'h294 == _way1_hit_T_1 ? cache_data_660 : _GEN_1683; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1685 = 10'h295 == _way1_hit_T_1 ? cache_data_661 : _GEN_1684; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1686 = 10'h296 == _way1_hit_T_1 ? cache_data_662 : _GEN_1685; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1687 = 10'h297 == _way1_hit_T_1 ? cache_data_663 : _GEN_1686; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1688 = 10'h298 == _way1_hit_T_1 ? cache_data_664 : _GEN_1687; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1689 = 10'h299 == _way1_hit_T_1 ? cache_data_665 : _GEN_1688; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1690 = 10'h29a == _way1_hit_T_1 ? cache_data_666 : _GEN_1689; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1691 = 10'h29b == _way1_hit_T_1 ? cache_data_667 : _GEN_1690; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1692 = 10'h29c == _way1_hit_T_1 ? cache_data_668 : _GEN_1691; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1693 = 10'h29d == _way1_hit_T_1 ? cache_data_669 : _GEN_1692; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1694 = 10'h29e == _way1_hit_T_1 ? cache_data_670 : _GEN_1693; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1695 = 10'h29f == _way1_hit_T_1 ? cache_data_671 : _GEN_1694; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1696 = 10'h2a0 == _way1_hit_T_1 ? cache_data_672 : _GEN_1695; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1697 = 10'h2a1 == _way1_hit_T_1 ? cache_data_673 : _GEN_1696; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1698 = 10'h2a2 == _way1_hit_T_1 ? cache_data_674 : _GEN_1697; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1699 = 10'h2a3 == _way1_hit_T_1 ? cache_data_675 : _GEN_1698; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1700 = 10'h2a4 == _way1_hit_T_1 ? cache_data_676 : _GEN_1699; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1701 = 10'h2a5 == _way1_hit_T_1 ? cache_data_677 : _GEN_1700; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1702 = 10'h2a6 == _way1_hit_T_1 ? cache_data_678 : _GEN_1701; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1703 = 10'h2a7 == _way1_hit_T_1 ? cache_data_679 : _GEN_1702; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1704 = 10'h2a8 == _way1_hit_T_1 ? cache_data_680 : _GEN_1703; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1705 = 10'h2a9 == _way1_hit_T_1 ? cache_data_681 : _GEN_1704; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1706 = 10'h2aa == _way1_hit_T_1 ? cache_data_682 : _GEN_1705; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1707 = 10'h2ab == _way1_hit_T_1 ? cache_data_683 : _GEN_1706; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1708 = 10'h2ac == _way1_hit_T_1 ? cache_data_684 : _GEN_1707; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1709 = 10'h2ad == _way1_hit_T_1 ? cache_data_685 : _GEN_1708; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1710 = 10'h2ae == _way1_hit_T_1 ? cache_data_686 : _GEN_1709; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1711 = 10'h2af == _way1_hit_T_1 ? cache_data_687 : _GEN_1710; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1712 = 10'h2b0 == _way1_hit_T_1 ? cache_data_688 : _GEN_1711; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1713 = 10'h2b1 == _way1_hit_T_1 ? cache_data_689 : _GEN_1712; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1714 = 10'h2b2 == _way1_hit_T_1 ? cache_data_690 : _GEN_1713; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1715 = 10'h2b3 == _way1_hit_T_1 ? cache_data_691 : _GEN_1714; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1716 = 10'h2b4 == _way1_hit_T_1 ? cache_data_692 : _GEN_1715; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1717 = 10'h2b5 == _way1_hit_T_1 ? cache_data_693 : _GEN_1716; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1718 = 10'h2b6 == _way1_hit_T_1 ? cache_data_694 : _GEN_1717; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1719 = 10'h2b7 == _way1_hit_T_1 ? cache_data_695 : _GEN_1718; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1720 = 10'h2b8 == _way1_hit_T_1 ? cache_data_696 : _GEN_1719; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1721 = 10'h2b9 == _way1_hit_T_1 ? cache_data_697 : _GEN_1720; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1722 = 10'h2ba == _way1_hit_T_1 ? cache_data_698 : _GEN_1721; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1723 = 10'h2bb == _way1_hit_T_1 ? cache_data_699 : _GEN_1722; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1724 = 10'h2bc == _way1_hit_T_1 ? cache_data_700 : _GEN_1723; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1725 = 10'h2bd == _way1_hit_T_1 ? cache_data_701 : _GEN_1724; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1726 = 10'h2be == _way1_hit_T_1 ? cache_data_702 : _GEN_1725; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1727 = 10'h2bf == _way1_hit_T_1 ? cache_data_703 : _GEN_1726; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1728 = 10'h2c0 == _way1_hit_T_1 ? cache_data_704 : _GEN_1727; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1729 = 10'h2c1 == _way1_hit_T_1 ? cache_data_705 : _GEN_1728; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1730 = 10'h2c2 == _way1_hit_T_1 ? cache_data_706 : _GEN_1729; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1731 = 10'h2c3 == _way1_hit_T_1 ? cache_data_707 : _GEN_1730; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1732 = 10'h2c4 == _way1_hit_T_1 ? cache_data_708 : _GEN_1731; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1733 = 10'h2c5 == _way1_hit_T_1 ? cache_data_709 : _GEN_1732; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1734 = 10'h2c6 == _way1_hit_T_1 ? cache_data_710 : _GEN_1733; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1735 = 10'h2c7 == _way1_hit_T_1 ? cache_data_711 : _GEN_1734; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1736 = 10'h2c8 == _way1_hit_T_1 ? cache_data_712 : _GEN_1735; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1737 = 10'h2c9 == _way1_hit_T_1 ? cache_data_713 : _GEN_1736; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1738 = 10'h2ca == _way1_hit_T_1 ? cache_data_714 : _GEN_1737; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1739 = 10'h2cb == _way1_hit_T_1 ? cache_data_715 : _GEN_1738; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1740 = 10'h2cc == _way1_hit_T_1 ? cache_data_716 : _GEN_1739; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1741 = 10'h2cd == _way1_hit_T_1 ? cache_data_717 : _GEN_1740; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1742 = 10'h2ce == _way1_hit_T_1 ? cache_data_718 : _GEN_1741; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1743 = 10'h2cf == _way1_hit_T_1 ? cache_data_719 : _GEN_1742; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1744 = 10'h2d0 == _way1_hit_T_1 ? cache_data_720 : _GEN_1743; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1745 = 10'h2d1 == _way1_hit_T_1 ? cache_data_721 : _GEN_1744; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1746 = 10'h2d2 == _way1_hit_T_1 ? cache_data_722 : _GEN_1745; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1747 = 10'h2d3 == _way1_hit_T_1 ? cache_data_723 : _GEN_1746; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1748 = 10'h2d4 == _way1_hit_T_1 ? cache_data_724 : _GEN_1747; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1749 = 10'h2d5 == _way1_hit_T_1 ? cache_data_725 : _GEN_1748; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1750 = 10'h2d6 == _way1_hit_T_1 ? cache_data_726 : _GEN_1749; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1751 = 10'h2d7 == _way1_hit_T_1 ? cache_data_727 : _GEN_1750; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1752 = 10'h2d8 == _way1_hit_T_1 ? cache_data_728 : _GEN_1751; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1753 = 10'h2d9 == _way1_hit_T_1 ? cache_data_729 : _GEN_1752; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1754 = 10'h2da == _way1_hit_T_1 ? cache_data_730 : _GEN_1753; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1755 = 10'h2db == _way1_hit_T_1 ? cache_data_731 : _GEN_1754; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1756 = 10'h2dc == _way1_hit_T_1 ? cache_data_732 : _GEN_1755; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1757 = 10'h2dd == _way1_hit_T_1 ? cache_data_733 : _GEN_1756; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1758 = 10'h2de == _way1_hit_T_1 ? cache_data_734 : _GEN_1757; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1759 = 10'h2df == _way1_hit_T_1 ? cache_data_735 : _GEN_1758; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1760 = 10'h2e0 == _way1_hit_T_1 ? cache_data_736 : _GEN_1759; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1761 = 10'h2e1 == _way1_hit_T_1 ? cache_data_737 : _GEN_1760; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1762 = 10'h2e2 == _way1_hit_T_1 ? cache_data_738 : _GEN_1761; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1763 = 10'h2e3 == _way1_hit_T_1 ? cache_data_739 : _GEN_1762; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1764 = 10'h2e4 == _way1_hit_T_1 ? cache_data_740 : _GEN_1763; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1765 = 10'h2e5 == _way1_hit_T_1 ? cache_data_741 : _GEN_1764; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1766 = 10'h2e6 == _way1_hit_T_1 ? cache_data_742 : _GEN_1765; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1767 = 10'h2e7 == _way1_hit_T_1 ? cache_data_743 : _GEN_1766; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1768 = 10'h2e8 == _way1_hit_T_1 ? cache_data_744 : _GEN_1767; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1769 = 10'h2e9 == _way1_hit_T_1 ? cache_data_745 : _GEN_1768; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1770 = 10'h2ea == _way1_hit_T_1 ? cache_data_746 : _GEN_1769; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1771 = 10'h2eb == _way1_hit_T_1 ? cache_data_747 : _GEN_1770; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1772 = 10'h2ec == _way1_hit_T_1 ? cache_data_748 : _GEN_1771; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1773 = 10'h2ed == _way1_hit_T_1 ? cache_data_749 : _GEN_1772; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1774 = 10'h2ee == _way1_hit_T_1 ? cache_data_750 : _GEN_1773; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1775 = 10'h2ef == _way1_hit_T_1 ? cache_data_751 : _GEN_1774; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1776 = 10'h2f0 == _way1_hit_T_1 ? cache_data_752 : _GEN_1775; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1777 = 10'h2f1 == _way1_hit_T_1 ? cache_data_753 : _GEN_1776; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1778 = 10'h2f2 == _way1_hit_T_1 ? cache_data_754 : _GEN_1777; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1779 = 10'h2f3 == _way1_hit_T_1 ? cache_data_755 : _GEN_1778; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1780 = 10'h2f4 == _way1_hit_T_1 ? cache_data_756 : _GEN_1779; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1781 = 10'h2f5 == _way1_hit_T_1 ? cache_data_757 : _GEN_1780; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1782 = 10'h2f6 == _way1_hit_T_1 ? cache_data_758 : _GEN_1781; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1783 = 10'h2f7 == _way1_hit_T_1 ? cache_data_759 : _GEN_1782; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1784 = 10'h2f8 == _way1_hit_T_1 ? cache_data_760 : _GEN_1783; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1785 = 10'h2f9 == _way1_hit_T_1 ? cache_data_761 : _GEN_1784; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1786 = 10'h2fa == _way1_hit_T_1 ? cache_data_762 : _GEN_1785; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1787 = 10'h2fb == _way1_hit_T_1 ? cache_data_763 : _GEN_1786; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1788 = 10'h2fc == _way1_hit_T_1 ? cache_data_764 : _GEN_1787; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1789 = 10'h2fd == _way1_hit_T_1 ? cache_data_765 : _GEN_1788; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1790 = 10'h2fe == _way1_hit_T_1 ? cache_data_766 : _GEN_1789; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1791 = 10'h2ff == _way1_hit_T_1 ? cache_data_767 : _GEN_1790; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1792 = 10'h300 == _way1_hit_T_1 ? cache_data_768 : _GEN_1791; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1793 = 10'h301 == _way1_hit_T_1 ? cache_data_769 : _GEN_1792; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1794 = 10'h302 == _way1_hit_T_1 ? cache_data_770 : _GEN_1793; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1795 = 10'h303 == _way1_hit_T_1 ? cache_data_771 : _GEN_1794; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1796 = 10'h304 == _way1_hit_T_1 ? cache_data_772 : _GEN_1795; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1797 = 10'h305 == _way1_hit_T_1 ? cache_data_773 : _GEN_1796; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1798 = 10'h306 == _way1_hit_T_1 ? cache_data_774 : _GEN_1797; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1799 = 10'h307 == _way1_hit_T_1 ? cache_data_775 : _GEN_1798; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1800 = 10'h308 == _way1_hit_T_1 ? cache_data_776 : _GEN_1799; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1801 = 10'h309 == _way1_hit_T_1 ? cache_data_777 : _GEN_1800; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1802 = 10'h30a == _way1_hit_T_1 ? cache_data_778 : _GEN_1801; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1803 = 10'h30b == _way1_hit_T_1 ? cache_data_779 : _GEN_1802; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1804 = 10'h30c == _way1_hit_T_1 ? cache_data_780 : _GEN_1803; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1805 = 10'h30d == _way1_hit_T_1 ? cache_data_781 : _GEN_1804; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1806 = 10'h30e == _way1_hit_T_1 ? cache_data_782 : _GEN_1805; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1807 = 10'h30f == _way1_hit_T_1 ? cache_data_783 : _GEN_1806; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1808 = 10'h310 == _way1_hit_T_1 ? cache_data_784 : _GEN_1807; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1809 = 10'h311 == _way1_hit_T_1 ? cache_data_785 : _GEN_1808; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1810 = 10'h312 == _way1_hit_T_1 ? cache_data_786 : _GEN_1809; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1811 = 10'h313 == _way1_hit_T_1 ? cache_data_787 : _GEN_1810; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1812 = 10'h314 == _way1_hit_T_1 ? cache_data_788 : _GEN_1811; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1813 = 10'h315 == _way1_hit_T_1 ? cache_data_789 : _GEN_1812; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1814 = 10'h316 == _way1_hit_T_1 ? cache_data_790 : _GEN_1813; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1815 = 10'h317 == _way1_hit_T_1 ? cache_data_791 : _GEN_1814; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1816 = 10'h318 == _way1_hit_T_1 ? cache_data_792 : _GEN_1815; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1817 = 10'h319 == _way1_hit_T_1 ? cache_data_793 : _GEN_1816; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1818 = 10'h31a == _way1_hit_T_1 ? cache_data_794 : _GEN_1817; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1819 = 10'h31b == _way1_hit_T_1 ? cache_data_795 : _GEN_1818; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1820 = 10'h31c == _way1_hit_T_1 ? cache_data_796 : _GEN_1819; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1821 = 10'h31d == _way1_hit_T_1 ? cache_data_797 : _GEN_1820; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1822 = 10'h31e == _way1_hit_T_1 ? cache_data_798 : _GEN_1821; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1823 = 10'h31f == _way1_hit_T_1 ? cache_data_799 : _GEN_1822; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1824 = 10'h320 == _way1_hit_T_1 ? cache_data_800 : _GEN_1823; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1825 = 10'h321 == _way1_hit_T_1 ? cache_data_801 : _GEN_1824; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1826 = 10'h322 == _way1_hit_T_1 ? cache_data_802 : _GEN_1825; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1827 = 10'h323 == _way1_hit_T_1 ? cache_data_803 : _GEN_1826; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1828 = 10'h324 == _way1_hit_T_1 ? cache_data_804 : _GEN_1827; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1829 = 10'h325 == _way1_hit_T_1 ? cache_data_805 : _GEN_1828; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1830 = 10'h326 == _way1_hit_T_1 ? cache_data_806 : _GEN_1829; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1831 = 10'h327 == _way1_hit_T_1 ? cache_data_807 : _GEN_1830; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1832 = 10'h328 == _way1_hit_T_1 ? cache_data_808 : _GEN_1831; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1833 = 10'h329 == _way1_hit_T_1 ? cache_data_809 : _GEN_1832; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1834 = 10'h32a == _way1_hit_T_1 ? cache_data_810 : _GEN_1833; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1835 = 10'h32b == _way1_hit_T_1 ? cache_data_811 : _GEN_1834; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1836 = 10'h32c == _way1_hit_T_1 ? cache_data_812 : _GEN_1835; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1837 = 10'h32d == _way1_hit_T_1 ? cache_data_813 : _GEN_1836; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1838 = 10'h32e == _way1_hit_T_1 ? cache_data_814 : _GEN_1837; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1839 = 10'h32f == _way1_hit_T_1 ? cache_data_815 : _GEN_1838; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1840 = 10'h330 == _way1_hit_T_1 ? cache_data_816 : _GEN_1839; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1841 = 10'h331 == _way1_hit_T_1 ? cache_data_817 : _GEN_1840; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1842 = 10'h332 == _way1_hit_T_1 ? cache_data_818 : _GEN_1841; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1843 = 10'h333 == _way1_hit_T_1 ? cache_data_819 : _GEN_1842; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1844 = 10'h334 == _way1_hit_T_1 ? cache_data_820 : _GEN_1843; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1845 = 10'h335 == _way1_hit_T_1 ? cache_data_821 : _GEN_1844; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1846 = 10'h336 == _way1_hit_T_1 ? cache_data_822 : _GEN_1845; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1847 = 10'h337 == _way1_hit_T_1 ? cache_data_823 : _GEN_1846; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1848 = 10'h338 == _way1_hit_T_1 ? cache_data_824 : _GEN_1847; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1849 = 10'h339 == _way1_hit_T_1 ? cache_data_825 : _GEN_1848; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1850 = 10'h33a == _way1_hit_T_1 ? cache_data_826 : _GEN_1849; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1851 = 10'h33b == _way1_hit_T_1 ? cache_data_827 : _GEN_1850; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1852 = 10'h33c == _way1_hit_T_1 ? cache_data_828 : _GEN_1851; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1853 = 10'h33d == _way1_hit_T_1 ? cache_data_829 : _GEN_1852; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1854 = 10'h33e == _way1_hit_T_1 ? cache_data_830 : _GEN_1853; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1855 = 10'h33f == _way1_hit_T_1 ? cache_data_831 : _GEN_1854; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1856 = 10'h340 == _way1_hit_T_1 ? cache_data_832 : _GEN_1855; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1857 = 10'h341 == _way1_hit_T_1 ? cache_data_833 : _GEN_1856; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1858 = 10'h342 == _way1_hit_T_1 ? cache_data_834 : _GEN_1857; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1859 = 10'h343 == _way1_hit_T_1 ? cache_data_835 : _GEN_1858; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1860 = 10'h344 == _way1_hit_T_1 ? cache_data_836 : _GEN_1859; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1861 = 10'h345 == _way1_hit_T_1 ? cache_data_837 : _GEN_1860; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1862 = 10'h346 == _way1_hit_T_1 ? cache_data_838 : _GEN_1861; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1863 = 10'h347 == _way1_hit_T_1 ? cache_data_839 : _GEN_1862; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1864 = 10'h348 == _way1_hit_T_1 ? cache_data_840 : _GEN_1863; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1865 = 10'h349 == _way1_hit_T_1 ? cache_data_841 : _GEN_1864; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1866 = 10'h34a == _way1_hit_T_1 ? cache_data_842 : _GEN_1865; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1867 = 10'h34b == _way1_hit_T_1 ? cache_data_843 : _GEN_1866; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1868 = 10'h34c == _way1_hit_T_1 ? cache_data_844 : _GEN_1867; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1869 = 10'h34d == _way1_hit_T_1 ? cache_data_845 : _GEN_1868; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1870 = 10'h34e == _way1_hit_T_1 ? cache_data_846 : _GEN_1869; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1871 = 10'h34f == _way1_hit_T_1 ? cache_data_847 : _GEN_1870; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1872 = 10'h350 == _way1_hit_T_1 ? cache_data_848 : _GEN_1871; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1873 = 10'h351 == _way1_hit_T_1 ? cache_data_849 : _GEN_1872; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1874 = 10'h352 == _way1_hit_T_1 ? cache_data_850 : _GEN_1873; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1875 = 10'h353 == _way1_hit_T_1 ? cache_data_851 : _GEN_1874; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1876 = 10'h354 == _way1_hit_T_1 ? cache_data_852 : _GEN_1875; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1877 = 10'h355 == _way1_hit_T_1 ? cache_data_853 : _GEN_1876; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1878 = 10'h356 == _way1_hit_T_1 ? cache_data_854 : _GEN_1877; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1879 = 10'h357 == _way1_hit_T_1 ? cache_data_855 : _GEN_1878; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1880 = 10'h358 == _way1_hit_T_1 ? cache_data_856 : _GEN_1879; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1881 = 10'h359 == _way1_hit_T_1 ? cache_data_857 : _GEN_1880; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1882 = 10'h35a == _way1_hit_T_1 ? cache_data_858 : _GEN_1881; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1883 = 10'h35b == _way1_hit_T_1 ? cache_data_859 : _GEN_1882; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1884 = 10'h35c == _way1_hit_T_1 ? cache_data_860 : _GEN_1883; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1885 = 10'h35d == _way1_hit_T_1 ? cache_data_861 : _GEN_1884; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1886 = 10'h35e == _way1_hit_T_1 ? cache_data_862 : _GEN_1885; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1887 = 10'h35f == _way1_hit_T_1 ? cache_data_863 : _GEN_1886; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1888 = 10'h360 == _way1_hit_T_1 ? cache_data_864 : _GEN_1887; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1889 = 10'h361 == _way1_hit_T_1 ? cache_data_865 : _GEN_1888; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1890 = 10'h362 == _way1_hit_T_1 ? cache_data_866 : _GEN_1889; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1891 = 10'h363 == _way1_hit_T_1 ? cache_data_867 : _GEN_1890; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1892 = 10'h364 == _way1_hit_T_1 ? cache_data_868 : _GEN_1891; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1893 = 10'h365 == _way1_hit_T_1 ? cache_data_869 : _GEN_1892; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1894 = 10'h366 == _way1_hit_T_1 ? cache_data_870 : _GEN_1893; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1895 = 10'h367 == _way1_hit_T_1 ? cache_data_871 : _GEN_1894; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1896 = 10'h368 == _way1_hit_T_1 ? cache_data_872 : _GEN_1895; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1897 = 10'h369 == _way1_hit_T_1 ? cache_data_873 : _GEN_1896; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1898 = 10'h36a == _way1_hit_T_1 ? cache_data_874 : _GEN_1897; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1899 = 10'h36b == _way1_hit_T_1 ? cache_data_875 : _GEN_1898; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1900 = 10'h36c == _way1_hit_T_1 ? cache_data_876 : _GEN_1899; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1901 = 10'h36d == _way1_hit_T_1 ? cache_data_877 : _GEN_1900; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1902 = 10'h36e == _way1_hit_T_1 ? cache_data_878 : _GEN_1901; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1903 = 10'h36f == _way1_hit_T_1 ? cache_data_879 : _GEN_1902; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1904 = 10'h370 == _way1_hit_T_1 ? cache_data_880 : _GEN_1903; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1905 = 10'h371 == _way1_hit_T_1 ? cache_data_881 : _GEN_1904; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1906 = 10'h372 == _way1_hit_T_1 ? cache_data_882 : _GEN_1905; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1907 = 10'h373 == _way1_hit_T_1 ? cache_data_883 : _GEN_1906; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1908 = 10'h374 == _way1_hit_T_1 ? cache_data_884 : _GEN_1907; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1909 = 10'h375 == _way1_hit_T_1 ? cache_data_885 : _GEN_1908; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1910 = 10'h376 == _way1_hit_T_1 ? cache_data_886 : _GEN_1909; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1911 = 10'h377 == _way1_hit_T_1 ? cache_data_887 : _GEN_1910; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1912 = 10'h378 == _way1_hit_T_1 ? cache_data_888 : _GEN_1911; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1913 = 10'h379 == _way1_hit_T_1 ? cache_data_889 : _GEN_1912; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1914 = 10'h37a == _way1_hit_T_1 ? cache_data_890 : _GEN_1913; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1915 = 10'h37b == _way1_hit_T_1 ? cache_data_891 : _GEN_1914; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1916 = 10'h37c == _way1_hit_T_1 ? cache_data_892 : _GEN_1915; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1917 = 10'h37d == _way1_hit_T_1 ? cache_data_893 : _GEN_1916; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1918 = 10'h37e == _way1_hit_T_1 ? cache_data_894 : _GEN_1917; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1919 = 10'h37f == _way1_hit_T_1 ? cache_data_895 : _GEN_1918; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1920 = 10'h380 == _way1_hit_T_1 ? cache_data_896 : _GEN_1919; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1921 = 10'h381 == _way1_hit_T_1 ? cache_data_897 : _GEN_1920; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1922 = 10'h382 == _way1_hit_T_1 ? cache_data_898 : _GEN_1921; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1923 = 10'h383 == _way1_hit_T_1 ? cache_data_899 : _GEN_1922; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1924 = 10'h384 == _way1_hit_T_1 ? cache_data_900 : _GEN_1923; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1925 = 10'h385 == _way1_hit_T_1 ? cache_data_901 : _GEN_1924; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1926 = 10'h386 == _way1_hit_T_1 ? cache_data_902 : _GEN_1925; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1927 = 10'h387 == _way1_hit_T_1 ? cache_data_903 : _GEN_1926; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1928 = 10'h388 == _way1_hit_T_1 ? cache_data_904 : _GEN_1927; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1929 = 10'h389 == _way1_hit_T_1 ? cache_data_905 : _GEN_1928; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1930 = 10'h38a == _way1_hit_T_1 ? cache_data_906 : _GEN_1929; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1931 = 10'h38b == _way1_hit_T_1 ? cache_data_907 : _GEN_1930; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1932 = 10'h38c == _way1_hit_T_1 ? cache_data_908 : _GEN_1931; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1933 = 10'h38d == _way1_hit_T_1 ? cache_data_909 : _GEN_1932; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1934 = 10'h38e == _way1_hit_T_1 ? cache_data_910 : _GEN_1933; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1935 = 10'h38f == _way1_hit_T_1 ? cache_data_911 : _GEN_1934; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1936 = 10'h390 == _way1_hit_T_1 ? cache_data_912 : _GEN_1935; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1937 = 10'h391 == _way1_hit_T_1 ? cache_data_913 : _GEN_1936; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1938 = 10'h392 == _way1_hit_T_1 ? cache_data_914 : _GEN_1937; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1939 = 10'h393 == _way1_hit_T_1 ? cache_data_915 : _GEN_1938; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1940 = 10'h394 == _way1_hit_T_1 ? cache_data_916 : _GEN_1939; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1941 = 10'h395 == _way1_hit_T_1 ? cache_data_917 : _GEN_1940; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1942 = 10'h396 == _way1_hit_T_1 ? cache_data_918 : _GEN_1941; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1943 = 10'h397 == _way1_hit_T_1 ? cache_data_919 : _GEN_1942; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1944 = 10'h398 == _way1_hit_T_1 ? cache_data_920 : _GEN_1943; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1945 = 10'h399 == _way1_hit_T_1 ? cache_data_921 : _GEN_1944; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1946 = 10'h39a == _way1_hit_T_1 ? cache_data_922 : _GEN_1945; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1947 = 10'h39b == _way1_hit_T_1 ? cache_data_923 : _GEN_1946; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1948 = 10'h39c == _way1_hit_T_1 ? cache_data_924 : _GEN_1947; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1949 = 10'h39d == _way1_hit_T_1 ? cache_data_925 : _GEN_1948; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1950 = 10'h39e == _way1_hit_T_1 ? cache_data_926 : _GEN_1949; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1951 = 10'h39f == _way1_hit_T_1 ? cache_data_927 : _GEN_1950; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1952 = 10'h3a0 == _way1_hit_T_1 ? cache_data_928 : _GEN_1951; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1953 = 10'h3a1 == _way1_hit_T_1 ? cache_data_929 : _GEN_1952; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1954 = 10'h3a2 == _way1_hit_T_1 ? cache_data_930 : _GEN_1953; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1955 = 10'h3a3 == _way1_hit_T_1 ? cache_data_931 : _GEN_1954; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1956 = 10'h3a4 == _way1_hit_T_1 ? cache_data_932 : _GEN_1955; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1957 = 10'h3a5 == _way1_hit_T_1 ? cache_data_933 : _GEN_1956; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1958 = 10'h3a6 == _way1_hit_T_1 ? cache_data_934 : _GEN_1957; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1959 = 10'h3a7 == _way1_hit_T_1 ? cache_data_935 : _GEN_1958; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1960 = 10'h3a8 == _way1_hit_T_1 ? cache_data_936 : _GEN_1959; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1961 = 10'h3a9 == _way1_hit_T_1 ? cache_data_937 : _GEN_1960; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1962 = 10'h3aa == _way1_hit_T_1 ? cache_data_938 : _GEN_1961; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1963 = 10'h3ab == _way1_hit_T_1 ? cache_data_939 : _GEN_1962; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1964 = 10'h3ac == _way1_hit_T_1 ? cache_data_940 : _GEN_1963; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1965 = 10'h3ad == _way1_hit_T_1 ? cache_data_941 : _GEN_1964; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1966 = 10'h3ae == _way1_hit_T_1 ? cache_data_942 : _GEN_1965; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1967 = 10'h3af == _way1_hit_T_1 ? cache_data_943 : _GEN_1966; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1968 = 10'h3b0 == _way1_hit_T_1 ? cache_data_944 : _GEN_1967; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1969 = 10'h3b1 == _way1_hit_T_1 ? cache_data_945 : _GEN_1968; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1970 = 10'h3b2 == _way1_hit_T_1 ? cache_data_946 : _GEN_1969; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1971 = 10'h3b3 == _way1_hit_T_1 ? cache_data_947 : _GEN_1970; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1972 = 10'h3b4 == _way1_hit_T_1 ? cache_data_948 : _GEN_1971; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1973 = 10'h3b5 == _way1_hit_T_1 ? cache_data_949 : _GEN_1972; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1974 = 10'h3b6 == _way1_hit_T_1 ? cache_data_950 : _GEN_1973; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1975 = 10'h3b7 == _way1_hit_T_1 ? cache_data_951 : _GEN_1974; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1976 = 10'h3b8 == _way1_hit_T_1 ? cache_data_952 : _GEN_1975; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1977 = 10'h3b9 == _way1_hit_T_1 ? cache_data_953 : _GEN_1976; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1978 = 10'h3ba == _way1_hit_T_1 ? cache_data_954 : _GEN_1977; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1979 = 10'h3bb == _way1_hit_T_1 ? cache_data_955 : _GEN_1978; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1980 = 10'h3bc == _way1_hit_T_1 ? cache_data_956 : _GEN_1979; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1981 = 10'h3bd == _way1_hit_T_1 ? cache_data_957 : _GEN_1980; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1982 = 10'h3be == _way1_hit_T_1 ? cache_data_958 : _GEN_1981; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1983 = 10'h3bf == _way1_hit_T_1 ? cache_data_959 : _GEN_1982; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1984 = 10'h3c0 == _way1_hit_T_1 ? cache_data_960 : _GEN_1983; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1985 = 10'h3c1 == _way1_hit_T_1 ? cache_data_961 : _GEN_1984; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1986 = 10'h3c2 == _way1_hit_T_1 ? cache_data_962 : _GEN_1985; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1987 = 10'h3c3 == _way1_hit_T_1 ? cache_data_963 : _GEN_1986; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1988 = 10'h3c4 == _way1_hit_T_1 ? cache_data_964 : _GEN_1987; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1989 = 10'h3c5 == _way1_hit_T_1 ? cache_data_965 : _GEN_1988; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1990 = 10'h3c6 == _way1_hit_T_1 ? cache_data_966 : _GEN_1989; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1991 = 10'h3c7 == _way1_hit_T_1 ? cache_data_967 : _GEN_1990; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1992 = 10'h3c8 == _way1_hit_T_1 ? cache_data_968 : _GEN_1991; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1993 = 10'h3c9 == _way1_hit_T_1 ? cache_data_969 : _GEN_1992; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1994 = 10'h3ca == _way1_hit_T_1 ? cache_data_970 : _GEN_1993; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1995 = 10'h3cb == _way1_hit_T_1 ? cache_data_971 : _GEN_1994; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1996 = 10'h3cc == _way1_hit_T_1 ? cache_data_972 : _GEN_1995; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1997 = 10'h3cd == _way1_hit_T_1 ? cache_data_973 : _GEN_1996; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1998 = 10'h3ce == _way1_hit_T_1 ? cache_data_974 : _GEN_1997; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_1999 = 10'h3cf == _way1_hit_T_1 ? cache_data_975 : _GEN_1998; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2000 = 10'h3d0 == _way1_hit_T_1 ? cache_data_976 : _GEN_1999; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2001 = 10'h3d1 == _way1_hit_T_1 ? cache_data_977 : _GEN_2000; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2002 = 10'h3d2 == _way1_hit_T_1 ? cache_data_978 : _GEN_2001; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2003 = 10'h3d3 == _way1_hit_T_1 ? cache_data_979 : _GEN_2002; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2004 = 10'h3d4 == _way1_hit_T_1 ? cache_data_980 : _GEN_2003; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2005 = 10'h3d5 == _way1_hit_T_1 ? cache_data_981 : _GEN_2004; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2006 = 10'h3d6 == _way1_hit_T_1 ? cache_data_982 : _GEN_2005; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2007 = 10'h3d7 == _way1_hit_T_1 ? cache_data_983 : _GEN_2006; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2008 = 10'h3d8 == _way1_hit_T_1 ? cache_data_984 : _GEN_2007; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2009 = 10'h3d9 == _way1_hit_T_1 ? cache_data_985 : _GEN_2008; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2010 = 10'h3da == _way1_hit_T_1 ? cache_data_986 : _GEN_2009; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2011 = 10'h3db == _way1_hit_T_1 ? cache_data_987 : _GEN_2010; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2012 = 10'h3dc == _way1_hit_T_1 ? cache_data_988 : _GEN_2011; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2013 = 10'h3dd == _way1_hit_T_1 ? cache_data_989 : _GEN_2012; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2014 = 10'h3de == _way1_hit_T_1 ? cache_data_990 : _GEN_2013; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2015 = 10'h3df == _way1_hit_T_1 ? cache_data_991 : _GEN_2014; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2016 = 10'h3e0 == _way1_hit_T_1 ? cache_data_992 : _GEN_2015; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2017 = 10'h3e1 == _way1_hit_T_1 ? cache_data_993 : _GEN_2016; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2018 = 10'h3e2 == _way1_hit_T_1 ? cache_data_994 : _GEN_2017; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2019 = 10'h3e3 == _way1_hit_T_1 ? cache_data_995 : _GEN_2018; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2020 = 10'h3e4 == _way1_hit_T_1 ? cache_data_996 : _GEN_2019; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2021 = 10'h3e5 == _way1_hit_T_1 ? cache_data_997 : _GEN_2020; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2022 = 10'h3e6 == _way1_hit_T_1 ? cache_data_998 : _GEN_2021; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2023 = 10'h3e7 == _way1_hit_T_1 ? cache_data_999 : _GEN_2022; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2024 = 10'h3e8 == _way1_hit_T_1 ? cache_data_1000 : _GEN_2023; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2025 = 10'h3e9 == _way1_hit_T_1 ? cache_data_1001 : _GEN_2024; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2026 = 10'h3ea == _way1_hit_T_1 ? cache_data_1002 : _GEN_2025; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2027 = 10'h3eb == _way1_hit_T_1 ? cache_data_1003 : _GEN_2026; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2028 = 10'h3ec == _way1_hit_T_1 ? cache_data_1004 : _GEN_2027; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2029 = 10'h3ed == _way1_hit_T_1 ? cache_data_1005 : _GEN_2028; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2030 = 10'h3ee == _way1_hit_T_1 ? cache_data_1006 : _GEN_2029; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2031 = 10'h3ef == _way1_hit_T_1 ? cache_data_1007 : _GEN_2030; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2032 = 10'h3f0 == _way1_hit_T_1 ? cache_data_1008 : _GEN_2031; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2033 = 10'h3f1 == _way1_hit_T_1 ? cache_data_1009 : _GEN_2032; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2034 = 10'h3f2 == _way1_hit_T_1 ? cache_data_1010 : _GEN_2033; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2035 = 10'h3f3 == _way1_hit_T_1 ? cache_data_1011 : _GEN_2034; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2036 = 10'h3f4 == _way1_hit_T_1 ? cache_data_1012 : _GEN_2035; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2037 = 10'h3f5 == _way1_hit_T_1 ? cache_data_1013 : _GEN_2036; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2038 = 10'h3f6 == _way1_hit_T_1 ? cache_data_1014 : _GEN_2037; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2039 = 10'h3f7 == _way1_hit_T_1 ? cache_data_1015 : _GEN_2038; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2040 = 10'h3f8 == _way1_hit_T_1 ? cache_data_1016 : _GEN_2039; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2041 = 10'h3f9 == _way1_hit_T_1 ? cache_data_1017 : _GEN_2040; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2042 = 10'h3fa == _way1_hit_T_1 ? cache_data_1018 : _GEN_2041; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2043 = 10'h3fb == _way1_hit_T_1 ? cache_data_1019 : _GEN_2042; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2044 = 10'h3fc == _way1_hit_T_1 ? cache_data_1020 : _GEN_2043; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2045 = 10'h3fd == _way1_hit_T_1 ? cache_data_1021 : _GEN_2044; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2046 = 10'h3fe == _way1_hit_T_1 ? cache_data_1022 : _GEN_2045; // @[icache.scala 49:{43,43}]
  wire [184:0] _GEN_2047 = 10'h3ff == _way1_hit_T_1 ? cache_data_1023 : _GEN_2046; // @[icache.scala 49:{43,43}]
  wire  way1_hit = _GEN_2047[184] & _GEN_2047[182:128] == cpu_tag; // @[icache.scala 49:58]
  wire  hit = way0_hit | way1_hit; // @[icache.scala 50:24]
  wire [1:0] _way_T_4 = {_GEN_1023[184],_GEN_2047[184]}; // @[Cat.scala 31:58]
  wire  _way_T_10 = 2'h3 == _way_T_4 | 2'h2 == _way_T_4; // @[Mux.scala 81:58]
  wire  way = ~hit & _way_T_10; // @[icache.scala 90:14 91:9]
  wire [9:0] _GEN_18450 = {{9'd0}, way}; // @[icache.scala 51:36]
  wire [9:0] _dirty_T_1 = cpu_index + _GEN_18450; // @[icache.scala 51:36]
  wire [184:0] _GEN_3073 = 10'h1 == _dirty_T_1 ? cache_data_1 : cache_data_0; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3074 = 10'h2 == _dirty_T_1 ? cache_data_2 : _GEN_3073; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3075 = 10'h3 == _dirty_T_1 ? cache_data_3 : _GEN_3074; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3076 = 10'h4 == _dirty_T_1 ? cache_data_4 : _GEN_3075; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3077 = 10'h5 == _dirty_T_1 ? cache_data_5 : _GEN_3076; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3078 = 10'h6 == _dirty_T_1 ? cache_data_6 : _GEN_3077; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3079 = 10'h7 == _dirty_T_1 ? cache_data_7 : _GEN_3078; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3080 = 10'h8 == _dirty_T_1 ? cache_data_8 : _GEN_3079; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3081 = 10'h9 == _dirty_T_1 ? cache_data_9 : _GEN_3080; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3082 = 10'ha == _dirty_T_1 ? cache_data_10 : _GEN_3081; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3083 = 10'hb == _dirty_T_1 ? cache_data_11 : _GEN_3082; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3084 = 10'hc == _dirty_T_1 ? cache_data_12 : _GEN_3083; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3085 = 10'hd == _dirty_T_1 ? cache_data_13 : _GEN_3084; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3086 = 10'he == _dirty_T_1 ? cache_data_14 : _GEN_3085; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3087 = 10'hf == _dirty_T_1 ? cache_data_15 : _GEN_3086; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3088 = 10'h10 == _dirty_T_1 ? cache_data_16 : _GEN_3087; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3089 = 10'h11 == _dirty_T_1 ? cache_data_17 : _GEN_3088; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3090 = 10'h12 == _dirty_T_1 ? cache_data_18 : _GEN_3089; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3091 = 10'h13 == _dirty_T_1 ? cache_data_19 : _GEN_3090; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3092 = 10'h14 == _dirty_T_1 ? cache_data_20 : _GEN_3091; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3093 = 10'h15 == _dirty_T_1 ? cache_data_21 : _GEN_3092; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3094 = 10'h16 == _dirty_T_1 ? cache_data_22 : _GEN_3093; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3095 = 10'h17 == _dirty_T_1 ? cache_data_23 : _GEN_3094; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3096 = 10'h18 == _dirty_T_1 ? cache_data_24 : _GEN_3095; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3097 = 10'h19 == _dirty_T_1 ? cache_data_25 : _GEN_3096; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3098 = 10'h1a == _dirty_T_1 ? cache_data_26 : _GEN_3097; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3099 = 10'h1b == _dirty_T_1 ? cache_data_27 : _GEN_3098; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3100 = 10'h1c == _dirty_T_1 ? cache_data_28 : _GEN_3099; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3101 = 10'h1d == _dirty_T_1 ? cache_data_29 : _GEN_3100; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3102 = 10'h1e == _dirty_T_1 ? cache_data_30 : _GEN_3101; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3103 = 10'h1f == _dirty_T_1 ? cache_data_31 : _GEN_3102; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3104 = 10'h20 == _dirty_T_1 ? cache_data_32 : _GEN_3103; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3105 = 10'h21 == _dirty_T_1 ? cache_data_33 : _GEN_3104; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3106 = 10'h22 == _dirty_T_1 ? cache_data_34 : _GEN_3105; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3107 = 10'h23 == _dirty_T_1 ? cache_data_35 : _GEN_3106; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3108 = 10'h24 == _dirty_T_1 ? cache_data_36 : _GEN_3107; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3109 = 10'h25 == _dirty_T_1 ? cache_data_37 : _GEN_3108; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3110 = 10'h26 == _dirty_T_1 ? cache_data_38 : _GEN_3109; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3111 = 10'h27 == _dirty_T_1 ? cache_data_39 : _GEN_3110; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3112 = 10'h28 == _dirty_T_1 ? cache_data_40 : _GEN_3111; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3113 = 10'h29 == _dirty_T_1 ? cache_data_41 : _GEN_3112; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3114 = 10'h2a == _dirty_T_1 ? cache_data_42 : _GEN_3113; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3115 = 10'h2b == _dirty_T_1 ? cache_data_43 : _GEN_3114; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3116 = 10'h2c == _dirty_T_1 ? cache_data_44 : _GEN_3115; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3117 = 10'h2d == _dirty_T_1 ? cache_data_45 : _GEN_3116; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3118 = 10'h2e == _dirty_T_1 ? cache_data_46 : _GEN_3117; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3119 = 10'h2f == _dirty_T_1 ? cache_data_47 : _GEN_3118; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3120 = 10'h30 == _dirty_T_1 ? cache_data_48 : _GEN_3119; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3121 = 10'h31 == _dirty_T_1 ? cache_data_49 : _GEN_3120; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3122 = 10'h32 == _dirty_T_1 ? cache_data_50 : _GEN_3121; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3123 = 10'h33 == _dirty_T_1 ? cache_data_51 : _GEN_3122; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3124 = 10'h34 == _dirty_T_1 ? cache_data_52 : _GEN_3123; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3125 = 10'h35 == _dirty_T_1 ? cache_data_53 : _GEN_3124; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3126 = 10'h36 == _dirty_T_1 ? cache_data_54 : _GEN_3125; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3127 = 10'h37 == _dirty_T_1 ? cache_data_55 : _GEN_3126; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3128 = 10'h38 == _dirty_T_1 ? cache_data_56 : _GEN_3127; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3129 = 10'h39 == _dirty_T_1 ? cache_data_57 : _GEN_3128; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3130 = 10'h3a == _dirty_T_1 ? cache_data_58 : _GEN_3129; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3131 = 10'h3b == _dirty_T_1 ? cache_data_59 : _GEN_3130; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3132 = 10'h3c == _dirty_T_1 ? cache_data_60 : _GEN_3131; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3133 = 10'h3d == _dirty_T_1 ? cache_data_61 : _GEN_3132; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3134 = 10'h3e == _dirty_T_1 ? cache_data_62 : _GEN_3133; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3135 = 10'h3f == _dirty_T_1 ? cache_data_63 : _GEN_3134; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3136 = 10'h40 == _dirty_T_1 ? cache_data_64 : _GEN_3135; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3137 = 10'h41 == _dirty_T_1 ? cache_data_65 : _GEN_3136; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3138 = 10'h42 == _dirty_T_1 ? cache_data_66 : _GEN_3137; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3139 = 10'h43 == _dirty_T_1 ? cache_data_67 : _GEN_3138; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3140 = 10'h44 == _dirty_T_1 ? cache_data_68 : _GEN_3139; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3141 = 10'h45 == _dirty_T_1 ? cache_data_69 : _GEN_3140; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3142 = 10'h46 == _dirty_T_1 ? cache_data_70 : _GEN_3141; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3143 = 10'h47 == _dirty_T_1 ? cache_data_71 : _GEN_3142; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3144 = 10'h48 == _dirty_T_1 ? cache_data_72 : _GEN_3143; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3145 = 10'h49 == _dirty_T_1 ? cache_data_73 : _GEN_3144; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3146 = 10'h4a == _dirty_T_1 ? cache_data_74 : _GEN_3145; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3147 = 10'h4b == _dirty_T_1 ? cache_data_75 : _GEN_3146; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3148 = 10'h4c == _dirty_T_1 ? cache_data_76 : _GEN_3147; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3149 = 10'h4d == _dirty_T_1 ? cache_data_77 : _GEN_3148; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3150 = 10'h4e == _dirty_T_1 ? cache_data_78 : _GEN_3149; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3151 = 10'h4f == _dirty_T_1 ? cache_data_79 : _GEN_3150; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3152 = 10'h50 == _dirty_T_1 ? cache_data_80 : _GEN_3151; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3153 = 10'h51 == _dirty_T_1 ? cache_data_81 : _GEN_3152; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3154 = 10'h52 == _dirty_T_1 ? cache_data_82 : _GEN_3153; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3155 = 10'h53 == _dirty_T_1 ? cache_data_83 : _GEN_3154; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3156 = 10'h54 == _dirty_T_1 ? cache_data_84 : _GEN_3155; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3157 = 10'h55 == _dirty_T_1 ? cache_data_85 : _GEN_3156; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3158 = 10'h56 == _dirty_T_1 ? cache_data_86 : _GEN_3157; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3159 = 10'h57 == _dirty_T_1 ? cache_data_87 : _GEN_3158; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3160 = 10'h58 == _dirty_T_1 ? cache_data_88 : _GEN_3159; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3161 = 10'h59 == _dirty_T_1 ? cache_data_89 : _GEN_3160; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3162 = 10'h5a == _dirty_T_1 ? cache_data_90 : _GEN_3161; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3163 = 10'h5b == _dirty_T_1 ? cache_data_91 : _GEN_3162; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3164 = 10'h5c == _dirty_T_1 ? cache_data_92 : _GEN_3163; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3165 = 10'h5d == _dirty_T_1 ? cache_data_93 : _GEN_3164; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3166 = 10'h5e == _dirty_T_1 ? cache_data_94 : _GEN_3165; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3167 = 10'h5f == _dirty_T_1 ? cache_data_95 : _GEN_3166; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3168 = 10'h60 == _dirty_T_1 ? cache_data_96 : _GEN_3167; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3169 = 10'h61 == _dirty_T_1 ? cache_data_97 : _GEN_3168; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3170 = 10'h62 == _dirty_T_1 ? cache_data_98 : _GEN_3169; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3171 = 10'h63 == _dirty_T_1 ? cache_data_99 : _GEN_3170; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3172 = 10'h64 == _dirty_T_1 ? cache_data_100 : _GEN_3171; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3173 = 10'h65 == _dirty_T_1 ? cache_data_101 : _GEN_3172; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3174 = 10'h66 == _dirty_T_1 ? cache_data_102 : _GEN_3173; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3175 = 10'h67 == _dirty_T_1 ? cache_data_103 : _GEN_3174; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3176 = 10'h68 == _dirty_T_1 ? cache_data_104 : _GEN_3175; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3177 = 10'h69 == _dirty_T_1 ? cache_data_105 : _GEN_3176; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3178 = 10'h6a == _dirty_T_1 ? cache_data_106 : _GEN_3177; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3179 = 10'h6b == _dirty_T_1 ? cache_data_107 : _GEN_3178; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3180 = 10'h6c == _dirty_T_1 ? cache_data_108 : _GEN_3179; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3181 = 10'h6d == _dirty_T_1 ? cache_data_109 : _GEN_3180; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3182 = 10'h6e == _dirty_T_1 ? cache_data_110 : _GEN_3181; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3183 = 10'h6f == _dirty_T_1 ? cache_data_111 : _GEN_3182; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3184 = 10'h70 == _dirty_T_1 ? cache_data_112 : _GEN_3183; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3185 = 10'h71 == _dirty_T_1 ? cache_data_113 : _GEN_3184; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3186 = 10'h72 == _dirty_T_1 ? cache_data_114 : _GEN_3185; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3187 = 10'h73 == _dirty_T_1 ? cache_data_115 : _GEN_3186; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3188 = 10'h74 == _dirty_T_1 ? cache_data_116 : _GEN_3187; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3189 = 10'h75 == _dirty_T_1 ? cache_data_117 : _GEN_3188; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3190 = 10'h76 == _dirty_T_1 ? cache_data_118 : _GEN_3189; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3191 = 10'h77 == _dirty_T_1 ? cache_data_119 : _GEN_3190; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3192 = 10'h78 == _dirty_T_1 ? cache_data_120 : _GEN_3191; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3193 = 10'h79 == _dirty_T_1 ? cache_data_121 : _GEN_3192; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3194 = 10'h7a == _dirty_T_1 ? cache_data_122 : _GEN_3193; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3195 = 10'h7b == _dirty_T_1 ? cache_data_123 : _GEN_3194; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3196 = 10'h7c == _dirty_T_1 ? cache_data_124 : _GEN_3195; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3197 = 10'h7d == _dirty_T_1 ? cache_data_125 : _GEN_3196; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3198 = 10'h7e == _dirty_T_1 ? cache_data_126 : _GEN_3197; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3199 = 10'h7f == _dirty_T_1 ? cache_data_127 : _GEN_3198; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3200 = 10'h80 == _dirty_T_1 ? cache_data_128 : _GEN_3199; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3201 = 10'h81 == _dirty_T_1 ? cache_data_129 : _GEN_3200; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3202 = 10'h82 == _dirty_T_1 ? cache_data_130 : _GEN_3201; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3203 = 10'h83 == _dirty_T_1 ? cache_data_131 : _GEN_3202; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3204 = 10'h84 == _dirty_T_1 ? cache_data_132 : _GEN_3203; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3205 = 10'h85 == _dirty_T_1 ? cache_data_133 : _GEN_3204; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3206 = 10'h86 == _dirty_T_1 ? cache_data_134 : _GEN_3205; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3207 = 10'h87 == _dirty_T_1 ? cache_data_135 : _GEN_3206; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3208 = 10'h88 == _dirty_T_1 ? cache_data_136 : _GEN_3207; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3209 = 10'h89 == _dirty_T_1 ? cache_data_137 : _GEN_3208; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3210 = 10'h8a == _dirty_T_1 ? cache_data_138 : _GEN_3209; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3211 = 10'h8b == _dirty_T_1 ? cache_data_139 : _GEN_3210; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3212 = 10'h8c == _dirty_T_1 ? cache_data_140 : _GEN_3211; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3213 = 10'h8d == _dirty_T_1 ? cache_data_141 : _GEN_3212; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3214 = 10'h8e == _dirty_T_1 ? cache_data_142 : _GEN_3213; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3215 = 10'h8f == _dirty_T_1 ? cache_data_143 : _GEN_3214; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3216 = 10'h90 == _dirty_T_1 ? cache_data_144 : _GEN_3215; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3217 = 10'h91 == _dirty_T_1 ? cache_data_145 : _GEN_3216; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3218 = 10'h92 == _dirty_T_1 ? cache_data_146 : _GEN_3217; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3219 = 10'h93 == _dirty_T_1 ? cache_data_147 : _GEN_3218; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3220 = 10'h94 == _dirty_T_1 ? cache_data_148 : _GEN_3219; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3221 = 10'h95 == _dirty_T_1 ? cache_data_149 : _GEN_3220; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3222 = 10'h96 == _dirty_T_1 ? cache_data_150 : _GEN_3221; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3223 = 10'h97 == _dirty_T_1 ? cache_data_151 : _GEN_3222; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3224 = 10'h98 == _dirty_T_1 ? cache_data_152 : _GEN_3223; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3225 = 10'h99 == _dirty_T_1 ? cache_data_153 : _GEN_3224; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3226 = 10'h9a == _dirty_T_1 ? cache_data_154 : _GEN_3225; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3227 = 10'h9b == _dirty_T_1 ? cache_data_155 : _GEN_3226; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3228 = 10'h9c == _dirty_T_1 ? cache_data_156 : _GEN_3227; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3229 = 10'h9d == _dirty_T_1 ? cache_data_157 : _GEN_3228; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3230 = 10'h9e == _dirty_T_1 ? cache_data_158 : _GEN_3229; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3231 = 10'h9f == _dirty_T_1 ? cache_data_159 : _GEN_3230; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3232 = 10'ha0 == _dirty_T_1 ? cache_data_160 : _GEN_3231; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3233 = 10'ha1 == _dirty_T_1 ? cache_data_161 : _GEN_3232; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3234 = 10'ha2 == _dirty_T_1 ? cache_data_162 : _GEN_3233; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3235 = 10'ha3 == _dirty_T_1 ? cache_data_163 : _GEN_3234; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3236 = 10'ha4 == _dirty_T_1 ? cache_data_164 : _GEN_3235; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3237 = 10'ha5 == _dirty_T_1 ? cache_data_165 : _GEN_3236; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3238 = 10'ha6 == _dirty_T_1 ? cache_data_166 : _GEN_3237; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3239 = 10'ha7 == _dirty_T_1 ? cache_data_167 : _GEN_3238; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3240 = 10'ha8 == _dirty_T_1 ? cache_data_168 : _GEN_3239; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3241 = 10'ha9 == _dirty_T_1 ? cache_data_169 : _GEN_3240; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3242 = 10'haa == _dirty_T_1 ? cache_data_170 : _GEN_3241; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3243 = 10'hab == _dirty_T_1 ? cache_data_171 : _GEN_3242; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3244 = 10'hac == _dirty_T_1 ? cache_data_172 : _GEN_3243; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3245 = 10'had == _dirty_T_1 ? cache_data_173 : _GEN_3244; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3246 = 10'hae == _dirty_T_1 ? cache_data_174 : _GEN_3245; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3247 = 10'haf == _dirty_T_1 ? cache_data_175 : _GEN_3246; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3248 = 10'hb0 == _dirty_T_1 ? cache_data_176 : _GEN_3247; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3249 = 10'hb1 == _dirty_T_1 ? cache_data_177 : _GEN_3248; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3250 = 10'hb2 == _dirty_T_1 ? cache_data_178 : _GEN_3249; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3251 = 10'hb3 == _dirty_T_1 ? cache_data_179 : _GEN_3250; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3252 = 10'hb4 == _dirty_T_1 ? cache_data_180 : _GEN_3251; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3253 = 10'hb5 == _dirty_T_1 ? cache_data_181 : _GEN_3252; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3254 = 10'hb6 == _dirty_T_1 ? cache_data_182 : _GEN_3253; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3255 = 10'hb7 == _dirty_T_1 ? cache_data_183 : _GEN_3254; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3256 = 10'hb8 == _dirty_T_1 ? cache_data_184 : _GEN_3255; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3257 = 10'hb9 == _dirty_T_1 ? cache_data_185 : _GEN_3256; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3258 = 10'hba == _dirty_T_1 ? cache_data_186 : _GEN_3257; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3259 = 10'hbb == _dirty_T_1 ? cache_data_187 : _GEN_3258; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3260 = 10'hbc == _dirty_T_1 ? cache_data_188 : _GEN_3259; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3261 = 10'hbd == _dirty_T_1 ? cache_data_189 : _GEN_3260; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3262 = 10'hbe == _dirty_T_1 ? cache_data_190 : _GEN_3261; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3263 = 10'hbf == _dirty_T_1 ? cache_data_191 : _GEN_3262; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3264 = 10'hc0 == _dirty_T_1 ? cache_data_192 : _GEN_3263; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3265 = 10'hc1 == _dirty_T_1 ? cache_data_193 : _GEN_3264; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3266 = 10'hc2 == _dirty_T_1 ? cache_data_194 : _GEN_3265; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3267 = 10'hc3 == _dirty_T_1 ? cache_data_195 : _GEN_3266; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3268 = 10'hc4 == _dirty_T_1 ? cache_data_196 : _GEN_3267; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3269 = 10'hc5 == _dirty_T_1 ? cache_data_197 : _GEN_3268; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3270 = 10'hc6 == _dirty_T_1 ? cache_data_198 : _GEN_3269; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3271 = 10'hc7 == _dirty_T_1 ? cache_data_199 : _GEN_3270; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3272 = 10'hc8 == _dirty_T_1 ? cache_data_200 : _GEN_3271; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3273 = 10'hc9 == _dirty_T_1 ? cache_data_201 : _GEN_3272; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3274 = 10'hca == _dirty_T_1 ? cache_data_202 : _GEN_3273; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3275 = 10'hcb == _dirty_T_1 ? cache_data_203 : _GEN_3274; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3276 = 10'hcc == _dirty_T_1 ? cache_data_204 : _GEN_3275; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3277 = 10'hcd == _dirty_T_1 ? cache_data_205 : _GEN_3276; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3278 = 10'hce == _dirty_T_1 ? cache_data_206 : _GEN_3277; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3279 = 10'hcf == _dirty_T_1 ? cache_data_207 : _GEN_3278; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3280 = 10'hd0 == _dirty_T_1 ? cache_data_208 : _GEN_3279; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3281 = 10'hd1 == _dirty_T_1 ? cache_data_209 : _GEN_3280; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3282 = 10'hd2 == _dirty_T_1 ? cache_data_210 : _GEN_3281; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3283 = 10'hd3 == _dirty_T_1 ? cache_data_211 : _GEN_3282; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3284 = 10'hd4 == _dirty_T_1 ? cache_data_212 : _GEN_3283; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3285 = 10'hd5 == _dirty_T_1 ? cache_data_213 : _GEN_3284; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3286 = 10'hd6 == _dirty_T_1 ? cache_data_214 : _GEN_3285; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3287 = 10'hd7 == _dirty_T_1 ? cache_data_215 : _GEN_3286; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3288 = 10'hd8 == _dirty_T_1 ? cache_data_216 : _GEN_3287; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3289 = 10'hd9 == _dirty_T_1 ? cache_data_217 : _GEN_3288; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3290 = 10'hda == _dirty_T_1 ? cache_data_218 : _GEN_3289; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3291 = 10'hdb == _dirty_T_1 ? cache_data_219 : _GEN_3290; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3292 = 10'hdc == _dirty_T_1 ? cache_data_220 : _GEN_3291; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3293 = 10'hdd == _dirty_T_1 ? cache_data_221 : _GEN_3292; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3294 = 10'hde == _dirty_T_1 ? cache_data_222 : _GEN_3293; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3295 = 10'hdf == _dirty_T_1 ? cache_data_223 : _GEN_3294; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3296 = 10'he0 == _dirty_T_1 ? cache_data_224 : _GEN_3295; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3297 = 10'he1 == _dirty_T_1 ? cache_data_225 : _GEN_3296; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3298 = 10'he2 == _dirty_T_1 ? cache_data_226 : _GEN_3297; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3299 = 10'he3 == _dirty_T_1 ? cache_data_227 : _GEN_3298; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3300 = 10'he4 == _dirty_T_1 ? cache_data_228 : _GEN_3299; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3301 = 10'he5 == _dirty_T_1 ? cache_data_229 : _GEN_3300; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3302 = 10'he6 == _dirty_T_1 ? cache_data_230 : _GEN_3301; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3303 = 10'he7 == _dirty_T_1 ? cache_data_231 : _GEN_3302; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3304 = 10'he8 == _dirty_T_1 ? cache_data_232 : _GEN_3303; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3305 = 10'he9 == _dirty_T_1 ? cache_data_233 : _GEN_3304; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3306 = 10'hea == _dirty_T_1 ? cache_data_234 : _GEN_3305; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3307 = 10'heb == _dirty_T_1 ? cache_data_235 : _GEN_3306; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3308 = 10'hec == _dirty_T_1 ? cache_data_236 : _GEN_3307; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3309 = 10'hed == _dirty_T_1 ? cache_data_237 : _GEN_3308; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3310 = 10'hee == _dirty_T_1 ? cache_data_238 : _GEN_3309; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3311 = 10'hef == _dirty_T_1 ? cache_data_239 : _GEN_3310; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3312 = 10'hf0 == _dirty_T_1 ? cache_data_240 : _GEN_3311; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3313 = 10'hf1 == _dirty_T_1 ? cache_data_241 : _GEN_3312; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3314 = 10'hf2 == _dirty_T_1 ? cache_data_242 : _GEN_3313; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3315 = 10'hf3 == _dirty_T_1 ? cache_data_243 : _GEN_3314; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3316 = 10'hf4 == _dirty_T_1 ? cache_data_244 : _GEN_3315; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3317 = 10'hf5 == _dirty_T_1 ? cache_data_245 : _GEN_3316; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3318 = 10'hf6 == _dirty_T_1 ? cache_data_246 : _GEN_3317; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3319 = 10'hf7 == _dirty_T_1 ? cache_data_247 : _GEN_3318; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3320 = 10'hf8 == _dirty_T_1 ? cache_data_248 : _GEN_3319; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3321 = 10'hf9 == _dirty_T_1 ? cache_data_249 : _GEN_3320; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3322 = 10'hfa == _dirty_T_1 ? cache_data_250 : _GEN_3321; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3323 = 10'hfb == _dirty_T_1 ? cache_data_251 : _GEN_3322; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3324 = 10'hfc == _dirty_T_1 ? cache_data_252 : _GEN_3323; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3325 = 10'hfd == _dirty_T_1 ? cache_data_253 : _GEN_3324; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3326 = 10'hfe == _dirty_T_1 ? cache_data_254 : _GEN_3325; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3327 = 10'hff == _dirty_T_1 ? cache_data_255 : _GEN_3326; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3328 = 10'h100 == _dirty_T_1 ? cache_data_256 : _GEN_3327; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3329 = 10'h101 == _dirty_T_1 ? cache_data_257 : _GEN_3328; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3330 = 10'h102 == _dirty_T_1 ? cache_data_258 : _GEN_3329; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3331 = 10'h103 == _dirty_T_1 ? cache_data_259 : _GEN_3330; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3332 = 10'h104 == _dirty_T_1 ? cache_data_260 : _GEN_3331; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3333 = 10'h105 == _dirty_T_1 ? cache_data_261 : _GEN_3332; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3334 = 10'h106 == _dirty_T_1 ? cache_data_262 : _GEN_3333; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3335 = 10'h107 == _dirty_T_1 ? cache_data_263 : _GEN_3334; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3336 = 10'h108 == _dirty_T_1 ? cache_data_264 : _GEN_3335; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3337 = 10'h109 == _dirty_T_1 ? cache_data_265 : _GEN_3336; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3338 = 10'h10a == _dirty_T_1 ? cache_data_266 : _GEN_3337; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3339 = 10'h10b == _dirty_T_1 ? cache_data_267 : _GEN_3338; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3340 = 10'h10c == _dirty_T_1 ? cache_data_268 : _GEN_3339; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3341 = 10'h10d == _dirty_T_1 ? cache_data_269 : _GEN_3340; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3342 = 10'h10e == _dirty_T_1 ? cache_data_270 : _GEN_3341; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3343 = 10'h10f == _dirty_T_1 ? cache_data_271 : _GEN_3342; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3344 = 10'h110 == _dirty_T_1 ? cache_data_272 : _GEN_3343; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3345 = 10'h111 == _dirty_T_1 ? cache_data_273 : _GEN_3344; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3346 = 10'h112 == _dirty_T_1 ? cache_data_274 : _GEN_3345; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3347 = 10'h113 == _dirty_T_1 ? cache_data_275 : _GEN_3346; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3348 = 10'h114 == _dirty_T_1 ? cache_data_276 : _GEN_3347; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3349 = 10'h115 == _dirty_T_1 ? cache_data_277 : _GEN_3348; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3350 = 10'h116 == _dirty_T_1 ? cache_data_278 : _GEN_3349; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3351 = 10'h117 == _dirty_T_1 ? cache_data_279 : _GEN_3350; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3352 = 10'h118 == _dirty_T_1 ? cache_data_280 : _GEN_3351; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3353 = 10'h119 == _dirty_T_1 ? cache_data_281 : _GEN_3352; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3354 = 10'h11a == _dirty_T_1 ? cache_data_282 : _GEN_3353; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3355 = 10'h11b == _dirty_T_1 ? cache_data_283 : _GEN_3354; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3356 = 10'h11c == _dirty_T_1 ? cache_data_284 : _GEN_3355; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3357 = 10'h11d == _dirty_T_1 ? cache_data_285 : _GEN_3356; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3358 = 10'h11e == _dirty_T_1 ? cache_data_286 : _GEN_3357; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3359 = 10'h11f == _dirty_T_1 ? cache_data_287 : _GEN_3358; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3360 = 10'h120 == _dirty_T_1 ? cache_data_288 : _GEN_3359; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3361 = 10'h121 == _dirty_T_1 ? cache_data_289 : _GEN_3360; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3362 = 10'h122 == _dirty_T_1 ? cache_data_290 : _GEN_3361; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3363 = 10'h123 == _dirty_T_1 ? cache_data_291 : _GEN_3362; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3364 = 10'h124 == _dirty_T_1 ? cache_data_292 : _GEN_3363; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3365 = 10'h125 == _dirty_T_1 ? cache_data_293 : _GEN_3364; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3366 = 10'h126 == _dirty_T_1 ? cache_data_294 : _GEN_3365; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3367 = 10'h127 == _dirty_T_1 ? cache_data_295 : _GEN_3366; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3368 = 10'h128 == _dirty_T_1 ? cache_data_296 : _GEN_3367; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3369 = 10'h129 == _dirty_T_1 ? cache_data_297 : _GEN_3368; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3370 = 10'h12a == _dirty_T_1 ? cache_data_298 : _GEN_3369; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3371 = 10'h12b == _dirty_T_1 ? cache_data_299 : _GEN_3370; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3372 = 10'h12c == _dirty_T_1 ? cache_data_300 : _GEN_3371; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3373 = 10'h12d == _dirty_T_1 ? cache_data_301 : _GEN_3372; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3374 = 10'h12e == _dirty_T_1 ? cache_data_302 : _GEN_3373; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3375 = 10'h12f == _dirty_T_1 ? cache_data_303 : _GEN_3374; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3376 = 10'h130 == _dirty_T_1 ? cache_data_304 : _GEN_3375; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3377 = 10'h131 == _dirty_T_1 ? cache_data_305 : _GEN_3376; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3378 = 10'h132 == _dirty_T_1 ? cache_data_306 : _GEN_3377; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3379 = 10'h133 == _dirty_T_1 ? cache_data_307 : _GEN_3378; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3380 = 10'h134 == _dirty_T_1 ? cache_data_308 : _GEN_3379; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3381 = 10'h135 == _dirty_T_1 ? cache_data_309 : _GEN_3380; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3382 = 10'h136 == _dirty_T_1 ? cache_data_310 : _GEN_3381; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3383 = 10'h137 == _dirty_T_1 ? cache_data_311 : _GEN_3382; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3384 = 10'h138 == _dirty_T_1 ? cache_data_312 : _GEN_3383; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3385 = 10'h139 == _dirty_T_1 ? cache_data_313 : _GEN_3384; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3386 = 10'h13a == _dirty_T_1 ? cache_data_314 : _GEN_3385; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3387 = 10'h13b == _dirty_T_1 ? cache_data_315 : _GEN_3386; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3388 = 10'h13c == _dirty_T_1 ? cache_data_316 : _GEN_3387; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3389 = 10'h13d == _dirty_T_1 ? cache_data_317 : _GEN_3388; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3390 = 10'h13e == _dirty_T_1 ? cache_data_318 : _GEN_3389; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3391 = 10'h13f == _dirty_T_1 ? cache_data_319 : _GEN_3390; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3392 = 10'h140 == _dirty_T_1 ? cache_data_320 : _GEN_3391; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3393 = 10'h141 == _dirty_T_1 ? cache_data_321 : _GEN_3392; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3394 = 10'h142 == _dirty_T_1 ? cache_data_322 : _GEN_3393; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3395 = 10'h143 == _dirty_T_1 ? cache_data_323 : _GEN_3394; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3396 = 10'h144 == _dirty_T_1 ? cache_data_324 : _GEN_3395; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3397 = 10'h145 == _dirty_T_1 ? cache_data_325 : _GEN_3396; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3398 = 10'h146 == _dirty_T_1 ? cache_data_326 : _GEN_3397; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3399 = 10'h147 == _dirty_T_1 ? cache_data_327 : _GEN_3398; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3400 = 10'h148 == _dirty_T_1 ? cache_data_328 : _GEN_3399; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3401 = 10'h149 == _dirty_T_1 ? cache_data_329 : _GEN_3400; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3402 = 10'h14a == _dirty_T_1 ? cache_data_330 : _GEN_3401; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3403 = 10'h14b == _dirty_T_1 ? cache_data_331 : _GEN_3402; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3404 = 10'h14c == _dirty_T_1 ? cache_data_332 : _GEN_3403; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3405 = 10'h14d == _dirty_T_1 ? cache_data_333 : _GEN_3404; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3406 = 10'h14e == _dirty_T_1 ? cache_data_334 : _GEN_3405; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3407 = 10'h14f == _dirty_T_1 ? cache_data_335 : _GEN_3406; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3408 = 10'h150 == _dirty_T_1 ? cache_data_336 : _GEN_3407; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3409 = 10'h151 == _dirty_T_1 ? cache_data_337 : _GEN_3408; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3410 = 10'h152 == _dirty_T_1 ? cache_data_338 : _GEN_3409; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3411 = 10'h153 == _dirty_T_1 ? cache_data_339 : _GEN_3410; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3412 = 10'h154 == _dirty_T_1 ? cache_data_340 : _GEN_3411; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3413 = 10'h155 == _dirty_T_1 ? cache_data_341 : _GEN_3412; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3414 = 10'h156 == _dirty_T_1 ? cache_data_342 : _GEN_3413; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3415 = 10'h157 == _dirty_T_1 ? cache_data_343 : _GEN_3414; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3416 = 10'h158 == _dirty_T_1 ? cache_data_344 : _GEN_3415; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3417 = 10'h159 == _dirty_T_1 ? cache_data_345 : _GEN_3416; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3418 = 10'h15a == _dirty_T_1 ? cache_data_346 : _GEN_3417; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3419 = 10'h15b == _dirty_T_1 ? cache_data_347 : _GEN_3418; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3420 = 10'h15c == _dirty_T_1 ? cache_data_348 : _GEN_3419; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3421 = 10'h15d == _dirty_T_1 ? cache_data_349 : _GEN_3420; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3422 = 10'h15e == _dirty_T_1 ? cache_data_350 : _GEN_3421; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3423 = 10'h15f == _dirty_T_1 ? cache_data_351 : _GEN_3422; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3424 = 10'h160 == _dirty_T_1 ? cache_data_352 : _GEN_3423; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3425 = 10'h161 == _dirty_T_1 ? cache_data_353 : _GEN_3424; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3426 = 10'h162 == _dirty_T_1 ? cache_data_354 : _GEN_3425; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3427 = 10'h163 == _dirty_T_1 ? cache_data_355 : _GEN_3426; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3428 = 10'h164 == _dirty_T_1 ? cache_data_356 : _GEN_3427; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3429 = 10'h165 == _dirty_T_1 ? cache_data_357 : _GEN_3428; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3430 = 10'h166 == _dirty_T_1 ? cache_data_358 : _GEN_3429; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3431 = 10'h167 == _dirty_T_1 ? cache_data_359 : _GEN_3430; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3432 = 10'h168 == _dirty_T_1 ? cache_data_360 : _GEN_3431; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3433 = 10'h169 == _dirty_T_1 ? cache_data_361 : _GEN_3432; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3434 = 10'h16a == _dirty_T_1 ? cache_data_362 : _GEN_3433; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3435 = 10'h16b == _dirty_T_1 ? cache_data_363 : _GEN_3434; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3436 = 10'h16c == _dirty_T_1 ? cache_data_364 : _GEN_3435; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3437 = 10'h16d == _dirty_T_1 ? cache_data_365 : _GEN_3436; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3438 = 10'h16e == _dirty_T_1 ? cache_data_366 : _GEN_3437; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3439 = 10'h16f == _dirty_T_1 ? cache_data_367 : _GEN_3438; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3440 = 10'h170 == _dirty_T_1 ? cache_data_368 : _GEN_3439; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3441 = 10'h171 == _dirty_T_1 ? cache_data_369 : _GEN_3440; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3442 = 10'h172 == _dirty_T_1 ? cache_data_370 : _GEN_3441; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3443 = 10'h173 == _dirty_T_1 ? cache_data_371 : _GEN_3442; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3444 = 10'h174 == _dirty_T_1 ? cache_data_372 : _GEN_3443; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3445 = 10'h175 == _dirty_T_1 ? cache_data_373 : _GEN_3444; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3446 = 10'h176 == _dirty_T_1 ? cache_data_374 : _GEN_3445; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3447 = 10'h177 == _dirty_T_1 ? cache_data_375 : _GEN_3446; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3448 = 10'h178 == _dirty_T_1 ? cache_data_376 : _GEN_3447; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3449 = 10'h179 == _dirty_T_1 ? cache_data_377 : _GEN_3448; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3450 = 10'h17a == _dirty_T_1 ? cache_data_378 : _GEN_3449; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3451 = 10'h17b == _dirty_T_1 ? cache_data_379 : _GEN_3450; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3452 = 10'h17c == _dirty_T_1 ? cache_data_380 : _GEN_3451; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3453 = 10'h17d == _dirty_T_1 ? cache_data_381 : _GEN_3452; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3454 = 10'h17e == _dirty_T_1 ? cache_data_382 : _GEN_3453; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3455 = 10'h17f == _dirty_T_1 ? cache_data_383 : _GEN_3454; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3456 = 10'h180 == _dirty_T_1 ? cache_data_384 : _GEN_3455; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3457 = 10'h181 == _dirty_T_1 ? cache_data_385 : _GEN_3456; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3458 = 10'h182 == _dirty_T_1 ? cache_data_386 : _GEN_3457; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3459 = 10'h183 == _dirty_T_1 ? cache_data_387 : _GEN_3458; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3460 = 10'h184 == _dirty_T_1 ? cache_data_388 : _GEN_3459; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3461 = 10'h185 == _dirty_T_1 ? cache_data_389 : _GEN_3460; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3462 = 10'h186 == _dirty_T_1 ? cache_data_390 : _GEN_3461; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3463 = 10'h187 == _dirty_T_1 ? cache_data_391 : _GEN_3462; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3464 = 10'h188 == _dirty_T_1 ? cache_data_392 : _GEN_3463; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3465 = 10'h189 == _dirty_T_1 ? cache_data_393 : _GEN_3464; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3466 = 10'h18a == _dirty_T_1 ? cache_data_394 : _GEN_3465; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3467 = 10'h18b == _dirty_T_1 ? cache_data_395 : _GEN_3466; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3468 = 10'h18c == _dirty_T_1 ? cache_data_396 : _GEN_3467; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3469 = 10'h18d == _dirty_T_1 ? cache_data_397 : _GEN_3468; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3470 = 10'h18e == _dirty_T_1 ? cache_data_398 : _GEN_3469; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3471 = 10'h18f == _dirty_T_1 ? cache_data_399 : _GEN_3470; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3472 = 10'h190 == _dirty_T_1 ? cache_data_400 : _GEN_3471; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3473 = 10'h191 == _dirty_T_1 ? cache_data_401 : _GEN_3472; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3474 = 10'h192 == _dirty_T_1 ? cache_data_402 : _GEN_3473; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3475 = 10'h193 == _dirty_T_1 ? cache_data_403 : _GEN_3474; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3476 = 10'h194 == _dirty_T_1 ? cache_data_404 : _GEN_3475; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3477 = 10'h195 == _dirty_T_1 ? cache_data_405 : _GEN_3476; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3478 = 10'h196 == _dirty_T_1 ? cache_data_406 : _GEN_3477; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3479 = 10'h197 == _dirty_T_1 ? cache_data_407 : _GEN_3478; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3480 = 10'h198 == _dirty_T_1 ? cache_data_408 : _GEN_3479; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3481 = 10'h199 == _dirty_T_1 ? cache_data_409 : _GEN_3480; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3482 = 10'h19a == _dirty_T_1 ? cache_data_410 : _GEN_3481; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3483 = 10'h19b == _dirty_T_1 ? cache_data_411 : _GEN_3482; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3484 = 10'h19c == _dirty_T_1 ? cache_data_412 : _GEN_3483; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3485 = 10'h19d == _dirty_T_1 ? cache_data_413 : _GEN_3484; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3486 = 10'h19e == _dirty_T_1 ? cache_data_414 : _GEN_3485; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3487 = 10'h19f == _dirty_T_1 ? cache_data_415 : _GEN_3486; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3488 = 10'h1a0 == _dirty_T_1 ? cache_data_416 : _GEN_3487; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3489 = 10'h1a1 == _dirty_T_1 ? cache_data_417 : _GEN_3488; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3490 = 10'h1a2 == _dirty_T_1 ? cache_data_418 : _GEN_3489; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3491 = 10'h1a3 == _dirty_T_1 ? cache_data_419 : _GEN_3490; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3492 = 10'h1a4 == _dirty_T_1 ? cache_data_420 : _GEN_3491; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3493 = 10'h1a5 == _dirty_T_1 ? cache_data_421 : _GEN_3492; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3494 = 10'h1a6 == _dirty_T_1 ? cache_data_422 : _GEN_3493; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3495 = 10'h1a7 == _dirty_T_1 ? cache_data_423 : _GEN_3494; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3496 = 10'h1a8 == _dirty_T_1 ? cache_data_424 : _GEN_3495; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3497 = 10'h1a9 == _dirty_T_1 ? cache_data_425 : _GEN_3496; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3498 = 10'h1aa == _dirty_T_1 ? cache_data_426 : _GEN_3497; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3499 = 10'h1ab == _dirty_T_1 ? cache_data_427 : _GEN_3498; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3500 = 10'h1ac == _dirty_T_1 ? cache_data_428 : _GEN_3499; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3501 = 10'h1ad == _dirty_T_1 ? cache_data_429 : _GEN_3500; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3502 = 10'h1ae == _dirty_T_1 ? cache_data_430 : _GEN_3501; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3503 = 10'h1af == _dirty_T_1 ? cache_data_431 : _GEN_3502; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3504 = 10'h1b0 == _dirty_T_1 ? cache_data_432 : _GEN_3503; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3505 = 10'h1b1 == _dirty_T_1 ? cache_data_433 : _GEN_3504; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3506 = 10'h1b2 == _dirty_T_1 ? cache_data_434 : _GEN_3505; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3507 = 10'h1b3 == _dirty_T_1 ? cache_data_435 : _GEN_3506; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3508 = 10'h1b4 == _dirty_T_1 ? cache_data_436 : _GEN_3507; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3509 = 10'h1b5 == _dirty_T_1 ? cache_data_437 : _GEN_3508; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3510 = 10'h1b6 == _dirty_T_1 ? cache_data_438 : _GEN_3509; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3511 = 10'h1b7 == _dirty_T_1 ? cache_data_439 : _GEN_3510; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3512 = 10'h1b8 == _dirty_T_1 ? cache_data_440 : _GEN_3511; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3513 = 10'h1b9 == _dirty_T_1 ? cache_data_441 : _GEN_3512; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3514 = 10'h1ba == _dirty_T_1 ? cache_data_442 : _GEN_3513; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3515 = 10'h1bb == _dirty_T_1 ? cache_data_443 : _GEN_3514; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3516 = 10'h1bc == _dirty_T_1 ? cache_data_444 : _GEN_3515; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3517 = 10'h1bd == _dirty_T_1 ? cache_data_445 : _GEN_3516; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3518 = 10'h1be == _dirty_T_1 ? cache_data_446 : _GEN_3517; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3519 = 10'h1bf == _dirty_T_1 ? cache_data_447 : _GEN_3518; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3520 = 10'h1c0 == _dirty_T_1 ? cache_data_448 : _GEN_3519; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3521 = 10'h1c1 == _dirty_T_1 ? cache_data_449 : _GEN_3520; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3522 = 10'h1c2 == _dirty_T_1 ? cache_data_450 : _GEN_3521; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3523 = 10'h1c3 == _dirty_T_1 ? cache_data_451 : _GEN_3522; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3524 = 10'h1c4 == _dirty_T_1 ? cache_data_452 : _GEN_3523; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3525 = 10'h1c5 == _dirty_T_1 ? cache_data_453 : _GEN_3524; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3526 = 10'h1c6 == _dirty_T_1 ? cache_data_454 : _GEN_3525; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3527 = 10'h1c7 == _dirty_T_1 ? cache_data_455 : _GEN_3526; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3528 = 10'h1c8 == _dirty_T_1 ? cache_data_456 : _GEN_3527; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3529 = 10'h1c9 == _dirty_T_1 ? cache_data_457 : _GEN_3528; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3530 = 10'h1ca == _dirty_T_1 ? cache_data_458 : _GEN_3529; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3531 = 10'h1cb == _dirty_T_1 ? cache_data_459 : _GEN_3530; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3532 = 10'h1cc == _dirty_T_1 ? cache_data_460 : _GEN_3531; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3533 = 10'h1cd == _dirty_T_1 ? cache_data_461 : _GEN_3532; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3534 = 10'h1ce == _dirty_T_1 ? cache_data_462 : _GEN_3533; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3535 = 10'h1cf == _dirty_T_1 ? cache_data_463 : _GEN_3534; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3536 = 10'h1d0 == _dirty_T_1 ? cache_data_464 : _GEN_3535; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3537 = 10'h1d1 == _dirty_T_1 ? cache_data_465 : _GEN_3536; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3538 = 10'h1d2 == _dirty_T_1 ? cache_data_466 : _GEN_3537; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3539 = 10'h1d3 == _dirty_T_1 ? cache_data_467 : _GEN_3538; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3540 = 10'h1d4 == _dirty_T_1 ? cache_data_468 : _GEN_3539; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3541 = 10'h1d5 == _dirty_T_1 ? cache_data_469 : _GEN_3540; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3542 = 10'h1d6 == _dirty_T_1 ? cache_data_470 : _GEN_3541; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3543 = 10'h1d7 == _dirty_T_1 ? cache_data_471 : _GEN_3542; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3544 = 10'h1d8 == _dirty_T_1 ? cache_data_472 : _GEN_3543; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3545 = 10'h1d9 == _dirty_T_1 ? cache_data_473 : _GEN_3544; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3546 = 10'h1da == _dirty_T_1 ? cache_data_474 : _GEN_3545; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3547 = 10'h1db == _dirty_T_1 ? cache_data_475 : _GEN_3546; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3548 = 10'h1dc == _dirty_T_1 ? cache_data_476 : _GEN_3547; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3549 = 10'h1dd == _dirty_T_1 ? cache_data_477 : _GEN_3548; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3550 = 10'h1de == _dirty_T_1 ? cache_data_478 : _GEN_3549; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3551 = 10'h1df == _dirty_T_1 ? cache_data_479 : _GEN_3550; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3552 = 10'h1e0 == _dirty_T_1 ? cache_data_480 : _GEN_3551; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3553 = 10'h1e1 == _dirty_T_1 ? cache_data_481 : _GEN_3552; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3554 = 10'h1e2 == _dirty_T_1 ? cache_data_482 : _GEN_3553; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3555 = 10'h1e3 == _dirty_T_1 ? cache_data_483 : _GEN_3554; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3556 = 10'h1e4 == _dirty_T_1 ? cache_data_484 : _GEN_3555; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3557 = 10'h1e5 == _dirty_T_1 ? cache_data_485 : _GEN_3556; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3558 = 10'h1e6 == _dirty_T_1 ? cache_data_486 : _GEN_3557; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3559 = 10'h1e7 == _dirty_T_1 ? cache_data_487 : _GEN_3558; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3560 = 10'h1e8 == _dirty_T_1 ? cache_data_488 : _GEN_3559; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3561 = 10'h1e9 == _dirty_T_1 ? cache_data_489 : _GEN_3560; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3562 = 10'h1ea == _dirty_T_1 ? cache_data_490 : _GEN_3561; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3563 = 10'h1eb == _dirty_T_1 ? cache_data_491 : _GEN_3562; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3564 = 10'h1ec == _dirty_T_1 ? cache_data_492 : _GEN_3563; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3565 = 10'h1ed == _dirty_T_1 ? cache_data_493 : _GEN_3564; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3566 = 10'h1ee == _dirty_T_1 ? cache_data_494 : _GEN_3565; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3567 = 10'h1ef == _dirty_T_1 ? cache_data_495 : _GEN_3566; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3568 = 10'h1f0 == _dirty_T_1 ? cache_data_496 : _GEN_3567; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3569 = 10'h1f1 == _dirty_T_1 ? cache_data_497 : _GEN_3568; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3570 = 10'h1f2 == _dirty_T_1 ? cache_data_498 : _GEN_3569; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3571 = 10'h1f3 == _dirty_T_1 ? cache_data_499 : _GEN_3570; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3572 = 10'h1f4 == _dirty_T_1 ? cache_data_500 : _GEN_3571; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3573 = 10'h1f5 == _dirty_T_1 ? cache_data_501 : _GEN_3572; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3574 = 10'h1f6 == _dirty_T_1 ? cache_data_502 : _GEN_3573; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3575 = 10'h1f7 == _dirty_T_1 ? cache_data_503 : _GEN_3574; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3576 = 10'h1f8 == _dirty_T_1 ? cache_data_504 : _GEN_3575; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3577 = 10'h1f9 == _dirty_T_1 ? cache_data_505 : _GEN_3576; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3578 = 10'h1fa == _dirty_T_1 ? cache_data_506 : _GEN_3577; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3579 = 10'h1fb == _dirty_T_1 ? cache_data_507 : _GEN_3578; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3580 = 10'h1fc == _dirty_T_1 ? cache_data_508 : _GEN_3579; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3581 = 10'h1fd == _dirty_T_1 ? cache_data_509 : _GEN_3580; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3582 = 10'h1fe == _dirty_T_1 ? cache_data_510 : _GEN_3581; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3583 = 10'h1ff == _dirty_T_1 ? cache_data_511 : _GEN_3582; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3584 = 10'h200 == _dirty_T_1 ? cache_data_512 : _GEN_3583; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3585 = 10'h201 == _dirty_T_1 ? cache_data_513 : _GEN_3584; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3586 = 10'h202 == _dirty_T_1 ? cache_data_514 : _GEN_3585; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3587 = 10'h203 == _dirty_T_1 ? cache_data_515 : _GEN_3586; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3588 = 10'h204 == _dirty_T_1 ? cache_data_516 : _GEN_3587; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3589 = 10'h205 == _dirty_T_1 ? cache_data_517 : _GEN_3588; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3590 = 10'h206 == _dirty_T_1 ? cache_data_518 : _GEN_3589; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3591 = 10'h207 == _dirty_T_1 ? cache_data_519 : _GEN_3590; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3592 = 10'h208 == _dirty_T_1 ? cache_data_520 : _GEN_3591; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3593 = 10'h209 == _dirty_T_1 ? cache_data_521 : _GEN_3592; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3594 = 10'h20a == _dirty_T_1 ? cache_data_522 : _GEN_3593; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3595 = 10'h20b == _dirty_T_1 ? cache_data_523 : _GEN_3594; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3596 = 10'h20c == _dirty_T_1 ? cache_data_524 : _GEN_3595; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3597 = 10'h20d == _dirty_T_1 ? cache_data_525 : _GEN_3596; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3598 = 10'h20e == _dirty_T_1 ? cache_data_526 : _GEN_3597; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3599 = 10'h20f == _dirty_T_1 ? cache_data_527 : _GEN_3598; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3600 = 10'h210 == _dirty_T_1 ? cache_data_528 : _GEN_3599; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3601 = 10'h211 == _dirty_T_1 ? cache_data_529 : _GEN_3600; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3602 = 10'h212 == _dirty_T_1 ? cache_data_530 : _GEN_3601; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3603 = 10'h213 == _dirty_T_1 ? cache_data_531 : _GEN_3602; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3604 = 10'h214 == _dirty_T_1 ? cache_data_532 : _GEN_3603; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3605 = 10'h215 == _dirty_T_1 ? cache_data_533 : _GEN_3604; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3606 = 10'h216 == _dirty_T_1 ? cache_data_534 : _GEN_3605; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3607 = 10'h217 == _dirty_T_1 ? cache_data_535 : _GEN_3606; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3608 = 10'h218 == _dirty_T_1 ? cache_data_536 : _GEN_3607; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3609 = 10'h219 == _dirty_T_1 ? cache_data_537 : _GEN_3608; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3610 = 10'h21a == _dirty_T_1 ? cache_data_538 : _GEN_3609; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3611 = 10'h21b == _dirty_T_1 ? cache_data_539 : _GEN_3610; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3612 = 10'h21c == _dirty_T_1 ? cache_data_540 : _GEN_3611; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3613 = 10'h21d == _dirty_T_1 ? cache_data_541 : _GEN_3612; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3614 = 10'h21e == _dirty_T_1 ? cache_data_542 : _GEN_3613; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3615 = 10'h21f == _dirty_T_1 ? cache_data_543 : _GEN_3614; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3616 = 10'h220 == _dirty_T_1 ? cache_data_544 : _GEN_3615; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3617 = 10'h221 == _dirty_T_1 ? cache_data_545 : _GEN_3616; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3618 = 10'h222 == _dirty_T_1 ? cache_data_546 : _GEN_3617; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3619 = 10'h223 == _dirty_T_1 ? cache_data_547 : _GEN_3618; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3620 = 10'h224 == _dirty_T_1 ? cache_data_548 : _GEN_3619; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3621 = 10'h225 == _dirty_T_1 ? cache_data_549 : _GEN_3620; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3622 = 10'h226 == _dirty_T_1 ? cache_data_550 : _GEN_3621; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3623 = 10'h227 == _dirty_T_1 ? cache_data_551 : _GEN_3622; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3624 = 10'h228 == _dirty_T_1 ? cache_data_552 : _GEN_3623; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3625 = 10'h229 == _dirty_T_1 ? cache_data_553 : _GEN_3624; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3626 = 10'h22a == _dirty_T_1 ? cache_data_554 : _GEN_3625; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3627 = 10'h22b == _dirty_T_1 ? cache_data_555 : _GEN_3626; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3628 = 10'h22c == _dirty_T_1 ? cache_data_556 : _GEN_3627; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3629 = 10'h22d == _dirty_T_1 ? cache_data_557 : _GEN_3628; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3630 = 10'h22e == _dirty_T_1 ? cache_data_558 : _GEN_3629; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3631 = 10'h22f == _dirty_T_1 ? cache_data_559 : _GEN_3630; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3632 = 10'h230 == _dirty_T_1 ? cache_data_560 : _GEN_3631; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3633 = 10'h231 == _dirty_T_1 ? cache_data_561 : _GEN_3632; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3634 = 10'h232 == _dirty_T_1 ? cache_data_562 : _GEN_3633; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3635 = 10'h233 == _dirty_T_1 ? cache_data_563 : _GEN_3634; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3636 = 10'h234 == _dirty_T_1 ? cache_data_564 : _GEN_3635; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3637 = 10'h235 == _dirty_T_1 ? cache_data_565 : _GEN_3636; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3638 = 10'h236 == _dirty_T_1 ? cache_data_566 : _GEN_3637; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3639 = 10'h237 == _dirty_T_1 ? cache_data_567 : _GEN_3638; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3640 = 10'h238 == _dirty_T_1 ? cache_data_568 : _GEN_3639; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3641 = 10'h239 == _dirty_T_1 ? cache_data_569 : _GEN_3640; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3642 = 10'h23a == _dirty_T_1 ? cache_data_570 : _GEN_3641; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3643 = 10'h23b == _dirty_T_1 ? cache_data_571 : _GEN_3642; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3644 = 10'h23c == _dirty_T_1 ? cache_data_572 : _GEN_3643; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3645 = 10'h23d == _dirty_T_1 ? cache_data_573 : _GEN_3644; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3646 = 10'h23e == _dirty_T_1 ? cache_data_574 : _GEN_3645; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3647 = 10'h23f == _dirty_T_1 ? cache_data_575 : _GEN_3646; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3648 = 10'h240 == _dirty_T_1 ? cache_data_576 : _GEN_3647; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3649 = 10'h241 == _dirty_T_1 ? cache_data_577 : _GEN_3648; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3650 = 10'h242 == _dirty_T_1 ? cache_data_578 : _GEN_3649; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3651 = 10'h243 == _dirty_T_1 ? cache_data_579 : _GEN_3650; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3652 = 10'h244 == _dirty_T_1 ? cache_data_580 : _GEN_3651; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3653 = 10'h245 == _dirty_T_1 ? cache_data_581 : _GEN_3652; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3654 = 10'h246 == _dirty_T_1 ? cache_data_582 : _GEN_3653; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3655 = 10'h247 == _dirty_T_1 ? cache_data_583 : _GEN_3654; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3656 = 10'h248 == _dirty_T_1 ? cache_data_584 : _GEN_3655; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3657 = 10'h249 == _dirty_T_1 ? cache_data_585 : _GEN_3656; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3658 = 10'h24a == _dirty_T_1 ? cache_data_586 : _GEN_3657; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3659 = 10'h24b == _dirty_T_1 ? cache_data_587 : _GEN_3658; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3660 = 10'h24c == _dirty_T_1 ? cache_data_588 : _GEN_3659; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3661 = 10'h24d == _dirty_T_1 ? cache_data_589 : _GEN_3660; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3662 = 10'h24e == _dirty_T_1 ? cache_data_590 : _GEN_3661; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3663 = 10'h24f == _dirty_T_1 ? cache_data_591 : _GEN_3662; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3664 = 10'h250 == _dirty_T_1 ? cache_data_592 : _GEN_3663; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3665 = 10'h251 == _dirty_T_1 ? cache_data_593 : _GEN_3664; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3666 = 10'h252 == _dirty_T_1 ? cache_data_594 : _GEN_3665; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3667 = 10'h253 == _dirty_T_1 ? cache_data_595 : _GEN_3666; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3668 = 10'h254 == _dirty_T_1 ? cache_data_596 : _GEN_3667; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3669 = 10'h255 == _dirty_T_1 ? cache_data_597 : _GEN_3668; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3670 = 10'h256 == _dirty_T_1 ? cache_data_598 : _GEN_3669; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3671 = 10'h257 == _dirty_T_1 ? cache_data_599 : _GEN_3670; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3672 = 10'h258 == _dirty_T_1 ? cache_data_600 : _GEN_3671; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3673 = 10'h259 == _dirty_T_1 ? cache_data_601 : _GEN_3672; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3674 = 10'h25a == _dirty_T_1 ? cache_data_602 : _GEN_3673; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3675 = 10'h25b == _dirty_T_1 ? cache_data_603 : _GEN_3674; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3676 = 10'h25c == _dirty_T_1 ? cache_data_604 : _GEN_3675; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3677 = 10'h25d == _dirty_T_1 ? cache_data_605 : _GEN_3676; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3678 = 10'h25e == _dirty_T_1 ? cache_data_606 : _GEN_3677; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3679 = 10'h25f == _dirty_T_1 ? cache_data_607 : _GEN_3678; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3680 = 10'h260 == _dirty_T_1 ? cache_data_608 : _GEN_3679; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3681 = 10'h261 == _dirty_T_1 ? cache_data_609 : _GEN_3680; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3682 = 10'h262 == _dirty_T_1 ? cache_data_610 : _GEN_3681; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3683 = 10'h263 == _dirty_T_1 ? cache_data_611 : _GEN_3682; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3684 = 10'h264 == _dirty_T_1 ? cache_data_612 : _GEN_3683; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3685 = 10'h265 == _dirty_T_1 ? cache_data_613 : _GEN_3684; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3686 = 10'h266 == _dirty_T_1 ? cache_data_614 : _GEN_3685; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3687 = 10'h267 == _dirty_T_1 ? cache_data_615 : _GEN_3686; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3688 = 10'h268 == _dirty_T_1 ? cache_data_616 : _GEN_3687; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3689 = 10'h269 == _dirty_T_1 ? cache_data_617 : _GEN_3688; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3690 = 10'h26a == _dirty_T_1 ? cache_data_618 : _GEN_3689; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3691 = 10'h26b == _dirty_T_1 ? cache_data_619 : _GEN_3690; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3692 = 10'h26c == _dirty_T_1 ? cache_data_620 : _GEN_3691; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3693 = 10'h26d == _dirty_T_1 ? cache_data_621 : _GEN_3692; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3694 = 10'h26e == _dirty_T_1 ? cache_data_622 : _GEN_3693; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3695 = 10'h26f == _dirty_T_1 ? cache_data_623 : _GEN_3694; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3696 = 10'h270 == _dirty_T_1 ? cache_data_624 : _GEN_3695; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3697 = 10'h271 == _dirty_T_1 ? cache_data_625 : _GEN_3696; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3698 = 10'h272 == _dirty_T_1 ? cache_data_626 : _GEN_3697; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3699 = 10'h273 == _dirty_T_1 ? cache_data_627 : _GEN_3698; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3700 = 10'h274 == _dirty_T_1 ? cache_data_628 : _GEN_3699; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3701 = 10'h275 == _dirty_T_1 ? cache_data_629 : _GEN_3700; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3702 = 10'h276 == _dirty_T_1 ? cache_data_630 : _GEN_3701; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3703 = 10'h277 == _dirty_T_1 ? cache_data_631 : _GEN_3702; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3704 = 10'h278 == _dirty_T_1 ? cache_data_632 : _GEN_3703; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3705 = 10'h279 == _dirty_T_1 ? cache_data_633 : _GEN_3704; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3706 = 10'h27a == _dirty_T_1 ? cache_data_634 : _GEN_3705; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3707 = 10'h27b == _dirty_T_1 ? cache_data_635 : _GEN_3706; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3708 = 10'h27c == _dirty_T_1 ? cache_data_636 : _GEN_3707; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3709 = 10'h27d == _dirty_T_1 ? cache_data_637 : _GEN_3708; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3710 = 10'h27e == _dirty_T_1 ? cache_data_638 : _GEN_3709; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3711 = 10'h27f == _dirty_T_1 ? cache_data_639 : _GEN_3710; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3712 = 10'h280 == _dirty_T_1 ? cache_data_640 : _GEN_3711; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3713 = 10'h281 == _dirty_T_1 ? cache_data_641 : _GEN_3712; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3714 = 10'h282 == _dirty_T_1 ? cache_data_642 : _GEN_3713; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3715 = 10'h283 == _dirty_T_1 ? cache_data_643 : _GEN_3714; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3716 = 10'h284 == _dirty_T_1 ? cache_data_644 : _GEN_3715; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3717 = 10'h285 == _dirty_T_1 ? cache_data_645 : _GEN_3716; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3718 = 10'h286 == _dirty_T_1 ? cache_data_646 : _GEN_3717; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3719 = 10'h287 == _dirty_T_1 ? cache_data_647 : _GEN_3718; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3720 = 10'h288 == _dirty_T_1 ? cache_data_648 : _GEN_3719; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3721 = 10'h289 == _dirty_T_1 ? cache_data_649 : _GEN_3720; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3722 = 10'h28a == _dirty_T_1 ? cache_data_650 : _GEN_3721; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3723 = 10'h28b == _dirty_T_1 ? cache_data_651 : _GEN_3722; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3724 = 10'h28c == _dirty_T_1 ? cache_data_652 : _GEN_3723; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3725 = 10'h28d == _dirty_T_1 ? cache_data_653 : _GEN_3724; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3726 = 10'h28e == _dirty_T_1 ? cache_data_654 : _GEN_3725; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3727 = 10'h28f == _dirty_T_1 ? cache_data_655 : _GEN_3726; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3728 = 10'h290 == _dirty_T_1 ? cache_data_656 : _GEN_3727; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3729 = 10'h291 == _dirty_T_1 ? cache_data_657 : _GEN_3728; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3730 = 10'h292 == _dirty_T_1 ? cache_data_658 : _GEN_3729; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3731 = 10'h293 == _dirty_T_1 ? cache_data_659 : _GEN_3730; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3732 = 10'h294 == _dirty_T_1 ? cache_data_660 : _GEN_3731; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3733 = 10'h295 == _dirty_T_1 ? cache_data_661 : _GEN_3732; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3734 = 10'h296 == _dirty_T_1 ? cache_data_662 : _GEN_3733; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3735 = 10'h297 == _dirty_T_1 ? cache_data_663 : _GEN_3734; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3736 = 10'h298 == _dirty_T_1 ? cache_data_664 : _GEN_3735; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3737 = 10'h299 == _dirty_T_1 ? cache_data_665 : _GEN_3736; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3738 = 10'h29a == _dirty_T_1 ? cache_data_666 : _GEN_3737; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3739 = 10'h29b == _dirty_T_1 ? cache_data_667 : _GEN_3738; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3740 = 10'h29c == _dirty_T_1 ? cache_data_668 : _GEN_3739; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3741 = 10'h29d == _dirty_T_1 ? cache_data_669 : _GEN_3740; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3742 = 10'h29e == _dirty_T_1 ? cache_data_670 : _GEN_3741; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3743 = 10'h29f == _dirty_T_1 ? cache_data_671 : _GEN_3742; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3744 = 10'h2a0 == _dirty_T_1 ? cache_data_672 : _GEN_3743; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3745 = 10'h2a1 == _dirty_T_1 ? cache_data_673 : _GEN_3744; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3746 = 10'h2a2 == _dirty_T_1 ? cache_data_674 : _GEN_3745; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3747 = 10'h2a3 == _dirty_T_1 ? cache_data_675 : _GEN_3746; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3748 = 10'h2a4 == _dirty_T_1 ? cache_data_676 : _GEN_3747; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3749 = 10'h2a5 == _dirty_T_1 ? cache_data_677 : _GEN_3748; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3750 = 10'h2a6 == _dirty_T_1 ? cache_data_678 : _GEN_3749; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3751 = 10'h2a7 == _dirty_T_1 ? cache_data_679 : _GEN_3750; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3752 = 10'h2a8 == _dirty_T_1 ? cache_data_680 : _GEN_3751; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3753 = 10'h2a9 == _dirty_T_1 ? cache_data_681 : _GEN_3752; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3754 = 10'h2aa == _dirty_T_1 ? cache_data_682 : _GEN_3753; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3755 = 10'h2ab == _dirty_T_1 ? cache_data_683 : _GEN_3754; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3756 = 10'h2ac == _dirty_T_1 ? cache_data_684 : _GEN_3755; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3757 = 10'h2ad == _dirty_T_1 ? cache_data_685 : _GEN_3756; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3758 = 10'h2ae == _dirty_T_1 ? cache_data_686 : _GEN_3757; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3759 = 10'h2af == _dirty_T_1 ? cache_data_687 : _GEN_3758; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3760 = 10'h2b0 == _dirty_T_1 ? cache_data_688 : _GEN_3759; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3761 = 10'h2b1 == _dirty_T_1 ? cache_data_689 : _GEN_3760; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3762 = 10'h2b2 == _dirty_T_1 ? cache_data_690 : _GEN_3761; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3763 = 10'h2b3 == _dirty_T_1 ? cache_data_691 : _GEN_3762; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3764 = 10'h2b4 == _dirty_T_1 ? cache_data_692 : _GEN_3763; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3765 = 10'h2b5 == _dirty_T_1 ? cache_data_693 : _GEN_3764; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3766 = 10'h2b6 == _dirty_T_1 ? cache_data_694 : _GEN_3765; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3767 = 10'h2b7 == _dirty_T_1 ? cache_data_695 : _GEN_3766; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3768 = 10'h2b8 == _dirty_T_1 ? cache_data_696 : _GEN_3767; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3769 = 10'h2b9 == _dirty_T_1 ? cache_data_697 : _GEN_3768; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3770 = 10'h2ba == _dirty_T_1 ? cache_data_698 : _GEN_3769; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3771 = 10'h2bb == _dirty_T_1 ? cache_data_699 : _GEN_3770; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3772 = 10'h2bc == _dirty_T_1 ? cache_data_700 : _GEN_3771; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3773 = 10'h2bd == _dirty_T_1 ? cache_data_701 : _GEN_3772; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3774 = 10'h2be == _dirty_T_1 ? cache_data_702 : _GEN_3773; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3775 = 10'h2bf == _dirty_T_1 ? cache_data_703 : _GEN_3774; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3776 = 10'h2c0 == _dirty_T_1 ? cache_data_704 : _GEN_3775; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3777 = 10'h2c1 == _dirty_T_1 ? cache_data_705 : _GEN_3776; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3778 = 10'h2c2 == _dirty_T_1 ? cache_data_706 : _GEN_3777; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3779 = 10'h2c3 == _dirty_T_1 ? cache_data_707 : _GEN_3778; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3780 = 10'h2c4 == _dirty_T_1 ? cache_data_708 : _GEN_3779; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3781 = 10'h2c5 == _dirty_T_1 ? cache_data_709 : _GEN_3780; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3782 = 10'h2c6 == _dirty_T_1 ? cache_data_710 : _GEN_3781; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3783 = 10'h2c7 == _dirty_T_1 ? cache_data_711 : _GEN_3782; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3784 = 10'h2c8 == _dirty_T_1 ? cache_data_712 : _GEN_3783; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3785 = 10'h2c9 == _dirty_T_1 ? cache_data_713 : _GEN_3784; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3786 = 10'h2ca == _dirty_T_1 ? cache_data_714 : _GEN_3785; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3787 = 10'h2cb == _dirty_T_1 ? cache_data_715 : _GEN_3786; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3788 = 10'h2cc == _dirty_T_1 ? cache_data_716 : _GEN_3787; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3789 = 10'h2cd == _dirty_T_1 ? cache_data_717 : _GEN_3788; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3790 = 10'h2ce == _dirty_T_1 ? cache_data_718 : _GEN_3789; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3791 = 10'h2cf == _dirty_T_1 ? cache_data_719 : _GEN_3790; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3792 = 10'h2d0 == _dirty_T_1 ? cache_data_720 : _GEN_3791; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3793 = 10'h2d1 == _dirty_T_1 ? cache_data_721 : _GEN_3792; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3794 = 10'h2d2 == _dirty_T_1 ? cache_data_722 : _GEN_3793; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3795 = 10'h2d3 == _dirty_T_1 ? cache_data_723 : _GEN_3794; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3796 = 10'h2d4 == _dirty_T_1 ? cache_data_724 : _GEN_3795; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3797 = 10'h2d5 == _dirty_T_1 ? cache_data_725 : _GEN_3796; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3798 = 10'h2d6 == _dirty_T_1 ? cache_data_726 : _GEN_3797; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3799 = 10'h2d7 == _dirty_T_1 ? cache_data_727 : _GEN_3798; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3800 = 10'h2d8 == _dirty_T_1 ? cache_data_728 : _GEN_3799; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3801 = 10'h2d9 == _dirty_T_1 ? cache_data_729 : _GEN_3800; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3802 = 10'h2da == _dirty_T_1 ? cache_data_730 : _GEN_3801; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3803 = 10'h2db == _dirty_T_1 ? cache_data_731 : _GEN_3802; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3804 = 10'h2dc == _dirty_T_1 ? cache_data_732 : _GEN_3803; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3805 = 10'h2dd == _dirty_T_1 ? cache_data_733 : _GEN_3804; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3806 = 10'h2de == _dirty_T_1 ? cache_data_734 : _GEN_3805; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3807 = 10'h2df == _dirty_T_1 ? cache_data_735 : _GEN_3806; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3808 = 10'h2e0 == _dirty_T_1 ? cache_data_736 : _GEN_3807; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3809 = 10'h2e1 == _dirty_T_1 ? cache_data_737 : _GEN_3808; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3810 = 10'h2e2 == _dirty_T_1 ? cache_data_738 : _GEN_3809; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3811 = 10'h2e3 == _dirty_T_1 ? cache_data_739 : _GEN_3810; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3812 = 10'h2e4 == _dirty_T_1 ? cache_data_740 : _GEN_3811; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3813 = 10'h2e5 == _dirty_T_1 ? cache_data_741 : _GEN_3812; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3814 = 10'h2e6 == _dirty_T_1 ? cache_data_742 : _GEN_3813; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3815 = 10'h2e7 == _dirty_T_1 ? cache_data_743 : _GEN_3814; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3816 = 10'h2e8 == _dirty_T_1 ? cache_data_744 : _GEN_3815; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3817 = 10'h2e9 == _dirty_T_1 ? cache_data_745 : _GEN_3816; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3818 = 10'h2ea == _dirty_T_1 ? cache_data_746 : _GEN_3817; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3819 = 10'h2eb == _dirty_T_1 ? cache_data_747 : _GEN_3818; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3820 = 10'h2ec == _dirty_T_1 ? cache_data_748 : _GEN_3819; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3821 = 10'h2ed == _dirty_T_1 ? cache_data_749 : _GEN_3820; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3822 = 10'h2ee == _dirty_T_1 ? cache_data_750 : _GEN_3821; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3823 = 10'h2ef == _dirty_T_1 ? cache_data_751 : _GEN_3822; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3824 = 10'h2f0 == _dirty_T_1 ? cache_data_752 : _GEN_3823; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3825 = 10'h2f1 == _dirty_T_1 ? cache_data_753 : _GEN_3824; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3826 = 10'h2f2 == _dirty_T_1 ? cache_data_754 : _GEN_3825; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3827 = 10'h2f3 == _dirty_T_1 ? cache_data_755 : _GEN_3826; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3828 = 10'h2f4 == _dirty_T_1 ? cache_data_756 : _GEN_3827; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3829 = 10'h2f5 == _dirty_T_1 ? cache_data_757 : _GEN_3828; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3830 = 10'h2f6 == _dirty_T_1 ? cache_data_758 : _GEN_3829; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3831 = 10'h2f7 == _dirty_T_1 ? cache_data_759 : _GEN_3830; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3832 = 10'h2f8 == _dirty_T_1 ? cache_data_760 : _GEN_3831; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3833 = 10'h2f9 == _dirty_T_1 ? cache_data_761 : _GEN_3832; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3834 = 10'h2fa == _dirty_T_1 ? cache_data_762 : _GEN_3833; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3835 = 10'h2fb == _dirty_T_1 ? cache_data_763 : _GEN_3834; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3836 = 10'h2fc == _dirty_T_1 ? cache_data_764 : _GEN_3835; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3837 = 10'h2fd == _dirty_T_1 ? cache_data_765 : _GEN_3836; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3838 = 10'h2fe == _dirty_T_1 ? cache_data_766 : _GEN_3837; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3839 = 10'h2ff == _dirty_T_1 ? cache_data_767 : _GEN_3838; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3840 = 10'h300 == _dirty_T_1 ? cache_data_768 : _GEN_3839; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3841 = 10'h301 == _dirty_T_1 ? cache_data_769 : _GEN_3840; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3842 = 10'h302 == _dirty_T_1 ? cache_data_770 : _GEN_3841; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3843 = 10'h303 == _dirty_T_1 ? cache_data_771 : _GEN_3842; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3844 = 10'h304 == _dirty_T_1 ? cache_data_772 : _GEN_3843; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3845 = 10'h305 == _dirty_T_1 ? cache_data_773 : _GEN_3844; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3846 = 10'h306 == _dirty_T_1 ? cache_data_774 : _GEN_3845; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3847 = 10'h307 == _dirty_T_1 ? cache_data_775 : _GEN_3846; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3848 = 10'h308 == _dirty_T_1 ? cache_data_776 : _GEN_3847; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3849 = 10'h309 == _dirty_T_1 ? cache_data_777 : _GEN_3848; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3850 = 10'h30a == _dirty_T_1 ? cache_data_778 : _GEN_3849; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3851 = 10'h30b == _dirty_T_1 ? cache_data_779 : _GEN_3850; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3852 = 10'h30c == _dirty_T_1 ? cache_data_780 : _GEN_3851; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3853 = 10'h30d == _dirty_T_1 ? cache_data_781 : _GEN_3852; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3854 = 10'h30e == _dirty_T_1 ? cache_data_782 : _GEN_3853; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3855 = 10'h30f == _dirty_T_1 ? cache_data_783 : _GEN_3854; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3856 = 10'h310 == _dirty_T_1 ? cache_data_784 : _GEN_3855; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3857 = 10'h311 == _dirty_T_1 ? cache_data_785 : _GEN_3856; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3858 = 10'h312 == _dirty_T_1 ? cache_data_786 : _GEN_3857; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3859 = 10'h313 == _dirty_T_1 ? cache_data_787 : _GEN_3858; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3860 = 10'h314 == _dirty_T_1 ? cache_data_788 : _GEN_3859; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3861 = 10'h315 == _dirty_T_1 ? cache_data_789 : _GEN_3860; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3862 = 10'h316 == _dirty_T_1 ? cache_data_790 : _GEN_3861; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3863 = 10'h317 == _dirty_T_1 ? cache_data_791 : _GEN_3862; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3864 = 10'h318 == _dirty_T_1 ? cache_data_792 : _GEN_3863; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3865 = 10'h319 == _dirty_T_1 ? cache_data_793 : _GEN_3864; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3866 = 10'h31a == _dirty_T_1 ? cache_data_794 : _GEN_3865; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3867 = 10'h31b == _dirty_T_1 ? cache_data_795 : _GEN_3866; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3868 = 10'h31c == _dirty_T_1 ? cache_data_796 : _GEN_3867; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3869 = 10'h31d == _dirty_T_1 ? cache_data_797 : _GEN_3868; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3870 = 10'h31e == _dirty_T_1 ? cache_data_798 : _GEN_3869; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3871 = 10'h31f == _dirty_T_1 ? cache_data_799 : _GEN_3870; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3872 = 10'h320 == _dirty_T_1 ? cache_data_800 : _GEN_3871; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3873 = 10'h321 == _dirty_T_1 ? cache_data_801 : _GEN_3872; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3874 = 10'h322 == _dirty_T_1 ? cache_data_802 : _GEN_3873; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3875 = 10'h323 == _dirty_T_1 ? cache_data_803 : _GEN_3874; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3876 = 10'h324 == _dirty_T_1 ? cache_data_804 : _GEN_3875; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3877 = 10'h325 == _dirty_T_1 ? cache_data_805 : _GEN_3876; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3878 = 10'h326 == _dirty_T_1 ? cache_data_806 : _GEN_3877; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3879 = 10'h327 == _dirty_T_1 ? cache_data_807 : _GEN_3878; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3880 = 10'h328 == _dirty_T_1 ? cache_data_808 : _GEN_3879; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3881 = 10'h329 == _dirty_T_1 ? cache_data_809 : _GEN_3880; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3882 = 10'h32a == _dirty_T_1 ? cache_data_810 : _GEN_3881; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3883 = 10'h32b == _dirty_T_1 ? cache_data_811 : _GEN_3882; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3884 = 10'h32c == _dirty_T_1 ? cache_data_812 : _GEN_3883; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3885 = 10'h32d == _dirty_T_1 ? cache_data_813 : _GEN_3884; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3886 = 10'h32e == _dirty_T_1 ? cache_data_814 : _GEN_3885; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3887 = 10'h32f == _dirty_T_1 ? cache_data_815 : _GEN_3886; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3888 = 10'h330 == _dirty_T_1 ? cache_data_816 : _GEN_3887; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3889 = 10'h331 == _dirty_T_1 ? cache_data_817 : _GEN_3888; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3890 = 10'h332 == _dirty_T_1 ? cache_data_818 : _GEN_3889; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3891 = 10'h333 == _dirty_T_1 ? cache_data_819 : _GEN_3890; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3892 = 10'h334 == _dirty_T_1 ? cache_data_820 : _GEN_3891; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3893 = 10'h335 == _dirty_T_1 ? cache_data_821 : _GEN_3892; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3894 = 10'h336 == _dirty_T_1 ? cache_data_822 : _GEN_3893; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3895 = 10'h337 == _dirty_T_1 ? cache_data_823 : _GEN_3894; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3896 = 10'h338 == _dirty_T_1 ? cache_data_824 : _GEN_3895; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3897 = 10'h339 == _dirty_T_1 ? cache_data_825 : _GEN_3896; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3898 = 10'h33a == _dirty_T_1 ? cache_data_826 : _GEN_3897; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3899 = 10'h33b == _dirty_T_1 ? cache_data_827 : _GEN_3898; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3900 = 10'h33c == _dirty_T_1 ? cache_data_828 : _GEN_3899; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3901 = 10'h33d == _dirty_T_1 ? cache_data_829 : _GEN_3900; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3902 = 10'h33e == _dirty_T_1 ? cache_data_830 : _GEN_3901; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3903 = 10'h33f == _dirty_T_1 ? cache_data_831 : _GEN_3902; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3904 = 10'h340 == _dirty_T_1 ? cache_data_832 : _GEN_3903; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3905 = 10'h341 == _dirty_T_1 ? cache_data_833 : _GEN_3904; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3906 = 10'h342 == _dirty_T_1 ? cache_data_834 : _GEN_3905; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3907 = 10'h343 == _dirty_T_1 ? cache_data_835 : _GEN_3906; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3908 = 10'h344 == _dirty_T_1 ? cache_data_836 : _GEN_3907; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3909 = 10'h345 == _dirty_T_1 ? cache_data_837 : _GEN_3908; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3910 = 10'h346 == _dirty_T_1 ? cache_data_838 : _GEN_3909; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3911 = 10'h347 == _dirty_T_1 ? cache_data_839 : _GEN_3910; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3912 = 10'h348 == _dirty_T_1 ? cache_data_840 : _GEN_3911; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3913 = 10'h349 == _dirty_T_1 ? cache_data_841 : _GEN_3912; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3914 = 10'h34a == _dirty_T_1 ? cache_data_842 : _GEN_3913; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3915 = 10'h34b == _dirty_T_1 ? cache_data_843 : _GEN_3914; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3916 = 10'h34c == _dirty_T_1 ? cache_data_844 : _GEN_3915; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3917 = 10'h34d == _dirty_T_1 ? cache_data_845 : _GEN_3916; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3918 = 10'h34e == _dirty_T_1 ? cache_data_846 : _GEN_3917; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3919 = 10'h34f == _dirty_T_1 ? cache_data_847 : _GEN_3918; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3920 = 10'h350 == _dirty_T_1 ? cache_data_848 : _GEN_3919; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3921 = 10'h351 == _dirty_T_1 ? cache_data_849 : _GEN_3920; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3922 = 10'h352 == _dirty_T_1 ? cache_data_850 : _GEN_3921; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3923 = 10'h353 == _dirty_T_1 ? cache_data_851 : _GEN_3922; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3924 = 10'h354 == _dirty_T_1 ? cache_data_852 : _GEN_3923; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3925 = 10'h355 == _dirty_T_1 ? cache_data_853 : _GEN_3924; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3926 = 10'h356 == _dirty_T_1 ? cache_data_854 : _GEN_3925; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3927 = 10'h357 == _dirty_T_1 ? cache_data_855 : _GEN_3926; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3928 = 10'h358 == _dirty_T_1 ? cache_data_856 : _GEN_3927; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3929 = 10'h359 == _dirty_T_1 ? cache_data_857 : _GEN_3928; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3930 = 10'h35a == _dirty_T_1 ? cache_data_858 : _GEN_3929; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3931 = 10'h35b == _dirty_T_1 ? cache_data_859 : _GEN_3930; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3932 = 10'h35c == _dirty_T_1 ? cache_data_860 : _GEN_3931; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3933 = 10'h35d == _dirty_T_1 ? cache_data_861 : _GEN_3932; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3934 = 10'h35e == _dirty_T_1 ? cache_data_862 : _GEN_3933; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3935 = 10'h35f == _dirty_T_1 ? cache_data_863 : _GEN_3934; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3936 = 10'h360 == _dirty_T_1 ? cache_data_864 : _GEN_3935; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3937 = 10'h361 == _dirty_T_1 ? cache_data_865 : _GEN_3936; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3938 = 10'h362 == _dirty_T_1 ? cache_data_866 : _GEN_3937; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3939 = 10'h363 == _dirty_T_1 ? cache_data_867 : _GEN_3938; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3940 = 10'h364 == _dirty_T_1 ? cache_data_868 : _GEN_3939; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3941 = 10'h365 == _dirty_T_1 ? cache_data_869 : _GEN_3940; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3942 = 10'h366 == _dirty_T_1 ? cache_data_870 : _GEN_3941; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3943 = 10'h367 == _dirty_T_1 ? cache_data_871 : _GEN_3942; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3944 = 10'h368 == _dirty_T_1 ? cache_data_872 : _GEN_3943; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3945 = 10'h369 == _dirty_T_1 ? cache_data_873 : _GEN_3944; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3946 = 10'h36a == _dirty_T_1 ? cache_data_874 : _GEN_3945; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3947 = 10'h36b == _dirty_T_1 ? cache_data_875 : _GEN_3946; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3948 = 10'h36c == _dirty_T_1 ? cache_data_876 : _GEN_3947; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3949 = 10'h36d == _dirty_T_1 ? cache_data_877 : _GEN_3948; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3950 = 10'h36e == _dirty_T_1 ? cache_data_878 : _GEN_3949; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3951 = 10'h36f == _dirty_T_1 ? cache_data_879 : _GEN_3950; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3952 = 10'h370 == _dirty_T_1 ? cache_data_880 : _GEN_3951; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3953 = 10'h371 == _dirty_T_1 ? cache_data_881 : _GEN_3952; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3954 = 10'h372 == _dirty_T_1 ? cache_data_882 : _GEN_3953; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3955 = 10'h373 == _dirty_T_1 ? cache_data_883 : _GEN_3954; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3956 = 10'h374 == _dirty_T_1 ? cache_data_884 : _GEN_3955; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3957 = 10'h375 == _dirty_T_1 ? cache_data_885 : _GEN_3956; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3958 = 10'h376 == _dirty_T_1 ? cache_data_886 : _GEN_3957; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3959 = 10'h377 == _dirty_T_1 ? cache_data_887 : _GEN_3958; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3960 = 10'h378 == _dirty_T_1 ? cache_data_888 : _GEN_3959; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3961 = 10'h379 == _dirty_T_1 ? cache_data_889 : _GEN_3960; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3962 = 10'h37a == _dirty_T_1 ? cache_data_890 : _GEN_3961; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3963 = 10'h37b == _dirty_T_1 ? cache_data_891 : _GEN_3962; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3964 = 10'h37c == _dirty_T_1 ? cache_data_892 : _GEN_3963; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3965 = 10'h37d == _dirty_T_1 ? cache_data_893 : _GEN_3964; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3966 = 10'h37e == _dirty_T_1 ? cache_data_894 : _GEN_3965; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3967 = 10'h37f == _dirty_T_1 ? cache_data_895 : _GEN_3966; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3968 = 10'h380 == _dirty_T_1 ? cache_data_896 : _GEN_3967; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3969 = 10'h381 == _dirty_T_1 ? cache_data_897 : _GEN_3968; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3970 = 10'h382 == _dirty_T_1 ? cache_data_898 : _GEN_3969; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3971 = 10'h383 == _dirty_T_1 ? cache_data_899 : _GEN_3970; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3972 = 10'h384 == _dirty_T_1 ? cache_data_900 : _GEN_3971; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3973 = 10'h385 == _dirty_T_1 ? cache_data_901 : _GEN_3972; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3974 = 10'h386 == _dirty_T_1 ? cache_data_902 : _GEN_3973; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3975 = 10'h387 == _dirty_T_1 ? cache_data_903 : _GEN_3974; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3976 = 10'h388 == _dirty_T_1 ? cache_data_904 : _GEN_3975; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3977 = 10'h389 == _dirty_T_1 ? cache_data_905 : _GEN_3976; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3978 = 10'h38a == _dirty_T_1 ? cache_data_906 : _GEN_3977; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3979 = 10'h38b == _dirty_T_1 ? cache_data_907 : _GEN_3978; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3980 = 10'h38c == _dirty_T_1 ? cache_data_908 : _GEN_3979; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3981 = 10'h38d == _dirty_T_1 ? cache_data_909 : _GEN_3980; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3982 = 10'h38e == _dirty_T_1 ? cache_data_910 : _GEN_3981; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3983 = 10'h38f == _dirty_T_1 ? cache_data_911 : _GEN_3982; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3984 = 10'h390 == _dirty_T_1 ? cache_data_912 : _GEN_3983; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3985 = 10'h391 == _dirty_T_1 ? cache_data_913 : _GEN_3984; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3986 = 10'h392 == _dirty_T_1 ? cache_data_914 : _GEN_3985; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3987 = 10'h393 == _dirty_T_1 ? cache_data_915 : _GEN_3986; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3988 = 10'h394 == _dirty_T_1 ? cache_data_916 : _GEN_3987; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3989 = 10'h395 == _dirty_T_1 ? cache_data_917 : _GEN_3988; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3990 = 10'h396 == _dirty_T_1 ? cache_data_918 : _GEN_3989; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3991 = 10'h397 == _dirty_T_1 ? cache_data_919 : _GEN_3990; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3992 = 10'h398 == _dirty_T_1 ? cache_data_920 : _GEN_3991; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3993 = 10'h399 == _dirty_T_1 ? cache_data_921 : _GEN_3992; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3994 = 10'h39a == _dirty_T_1 ? cache_data_922 : _GEN_3993; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3995 = 10'h39b == _dirty_T_1 ? cache_data_923 : _GEN_3994; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3996 = 10'h39c == _dirty_T_1 ? cache_data_924 : _GEN_3995; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3997 = 10'h39d == _dirty_T_1 ? cache_data_925 : _GEN_3996; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3998 = 10'h39e == _dirty_T_1 ? cache_data_926 : _GEN_3997; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_3999 = 10'h39f == _dirty_T_1 ? cache_data_927 : _GEN_3998; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4000 = 10'h3a0 == _dirty_T_1 ? cache_data_928 : _GEN_3999; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4001 = 10'h3a1 == _dirty_T_1 ? cache_data_929 : _GEN_4000; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4002 = 10'h3a2 == _dirty_T_1 ? cache_data_930 : _GEN_4001; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4003 = 10'h3a3 == _dirty_T_1 ? cache_data_931 : _GEN_4002; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4004 = 10'h3a4 == _dirty_T_1 ? cache_data_932 : _GEN_4003; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4005 = 10'h3a5 == _dirty_T_1 ? cache_data_933 : _GEN_4004; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4006 = 10'h3a6 == _dirty_T_1 ? cache_data_934 : _GEN_4005; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4007 = 10'h3a7 == _dirty_T_1 ? cache_data_935 : _GEN_4006; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4008 = 10'h3a8 == _dirty_T_1 ? cache_data_936 : _GEN_4007; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4009 = 10'h3a9 == _dirty_T_1 ? cache_data_937 : _GEN_4008; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4010 = 10'h3aa == _dirty_T_1 ? cache_data_938 : _GEN_4009; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4011 = 10'h3ab == _dirty_T_1 ? cache_data_939 : _GEN_4010; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4012 = 10'h3ac == _dirty_T_1 ? cache_data_940 : _GEN_4011; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4013 = 10'h3ad == _dirty_T_1 ? cache_data_941 : _GEN_4012; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4014 = 10'h3ae == _dirty_T_1 ? cache_data_942 : _GEN_4013; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4015 = 10'h3af == _dirty_T_1 ? cache_data_943 : _GEN_4014; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4016 = 10'h3b0 == _dirty_T_1 ? cache_data_944 : _GEN_4015; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4017 = 10'h3b1 == _dirty_T_1 ? cache_data_945 : _GEN_4016; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4018 = 10'h3b2 == _dirty_T_1 ? cache_data_946 : _GEN_4017; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4019 = 10'h3b3 == _dirty_T_1 ? cache_data_947 : _GEN_4018; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4020 = 10'h3b4 == _dirty_T_1 ? cache_data_948 : _GEN_4019; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4021 = 10'h3b5 == _dirty_T_1 ? cache_data_949 : _GEN_4020; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4022 = 10'h3b6 == _dirty_T_1 ? cache_data_950 : _GEN_4021; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4023 = 10'h3b7 == _dirty_T_1 ? cache_data_951 : _GEN_4022; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4024 = 10'h3b8 == _dirty_T_1 ? cache_data_952 : _GEN_4023; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4025 = 10'h3b9 == _dirty_T_1 ? cache_data_953 : _GEN_4024; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4026 = 10'h3ba == _dirty_T_1 ? cache_data_954 : _GEN_4025; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4027 = 10'h3bb == _dirty_T_1 ? cache_data_955 : _GEN_4026; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4028 = 10'h3bc == _dirty_T_1 ? cache_data_956 : _GEN_4027; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4029 = 10'h3bd == _dirty_T_1 ? cache_data_957 : _GEN_4028; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4030 = 10'h3be == _dirty_T_1 ? cache_data_958 : _GEN_4029; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4031 = 10'h3bf == _dirty_T_1 ? cache_data_959 : _GEN_4030; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4032 = 10'h3c0 == _dirty_T_1 ? cache_data_960 : _GEN_4031; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4033 = 10'h3c1 == _dirty_T_1 ? cache_data_961 : _GEN_4032; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4034 = 10'h3c2 == _dirty_T_1 ? cache_data_962 : _GEN_4033; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4035 = 10'h3c3 == _dirty_T_1 ? cache_data_963 : _GEN_4034; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4036 = 10'h3c4 == _dirty_T_1 ? cache_data_964 : _GEN_4035; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4037 = 10'h3c5 == _dirty_T_1 ? cache_data_965 : _GEN_4036; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4038 = 10'h3c6 == _dirty_T_1 ? cache_data_966 : _GEN_4037; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4039 = 10'h3c7 == _dirty_T_1 ? cache_data_967 : _GEN_4038; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4040 = 10'h3c8 == _dirty_T_1 ? cache_data_968 : _GEN_4039; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4041 = 10'h3c9 == _dirty_T_1 ? cache_data_969 : _GEN_4040; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4042 = 10'h3ca == _dirty_T_1 ? cache_data_970 : _GEN_4041; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4043 = 10'h3cb == _dirty_T_1 ? cache_data_971 : _GEN_4042; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4044 = 10'h3cc == _dirty_T_1 ? cache_data_972 : _GEN_4043; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4045 = 10'h3cd == _dirty_T_1 ? cache_data_973 : _GEN_4044; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4046 = 10'h3ce == _dirty_T_1 ? cache_data_974 : _GEN_4045; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4047 = 10'h3cf == _dirty_T_1 ? cache_data_975 : _GEN_4046; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4048 = 10'h3d0 == _dirty_T_1 ? cache_data_976 : _GEN_4047; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4049 = 10'h3d1 == _dirty_T_1 ? cache_data_977 : _GEN_4048; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4050 = 10'h3d2 == _dirty_T_1 ? cache_data_978 : _GEN_4049; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4051 = 10'h3d3 == _dirty_T_1 ? cache_data_979 : _GEN_4050; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4052 = 10'h3d4 == _dirty_T_1 ? cache_data_980 : _GEN_4051; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4053 = 10'h3d5 == _dirty_T_1 ? cache_data_981 : _GEN_4052; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4054 = 10'h3d6 == _dirty_T_1 ? cache_data_982 : _GEN_4053; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4055 = 10'h3d7 == _dirty_T_1 ? cache_data_983 : _GEN_4054; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4056 = 10'h3d8 == _dirty_T_1 ? cache_data_984 : _GEN_4055; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4057 = 10'h3d9 == _dirty_T_1 ? cache_data_985 : _GEN_4056; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4058 = 10'h3da == _dirty_T_1 ? cache_data_986 : _GEN_4057; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4059 = 10'h3db == _dirty_T_1 ? cache_data_987 : _GEN_4058; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4060 = 10'h3dc == _dirty_T_1 ? cache_data_988 : _GEN_4059; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4061 = 10'h3dd == _dirty_T_1 ? cache_data_989 : _GEN_4060; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4062 = 10'h3de == _dirty_T_1 ? cache_data_990 : _GEN_4061; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4063 = 10'h3df == _dirty_T_1 ? cache_data_991 : _GEN_4062; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4064 = 10'h3e0 == _dirty_T_1 ? cache_data_992 : _GEN_4063; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4065 = 10'h3e1 == _dirty_T_1 ? cache_data_993 : _GEN_4064; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4066 = 10'h3e2 == _dirty_T_1 ? cache_data_994 : _GEN_4065; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4067 = 10'h3e3 == _dirty_T_1 ? cache_data_995 : _GEN_4066; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4068 = 10'h3e4 == _dirty_T_1 ? cache_data_996 : _GEN_4067; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4069 = 10'h3e5 == _dirty_T_1 ? cache_data_997 : _GEN_4068; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4070 = 10'h3e6 == _dirty_T_1 ? cache_data_998 : _GEN_4069; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4071 = 10'h3e7 == _dirty_T_1 ? cache_data_999 : _GEN_4070; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4072 = 10'h3e8 == _dirty_T_1 ? cache_data_1000 : _GEN_4071; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4073 = 10'h3e9 == _dirty_T_1 ? cache_data_1001 : _GEN_4072; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4074 = 10'h3ea == _dirty_T_1 ? cache_data_1002 : _GEN_4073; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4075 = 10'h3eb == _dirty_T_1 ? cache_data_1003 : _GEN_4074; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4076 = 10'h3ec == _dirty_T_1 ? cache_data_1004 : _GEN_4075; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4077 = 10'h3ed == _dirty_T_1 ? cache_data_1005 : _GEN_4076; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4078 = 10'h3ee == _dirty_T_1 ? cache_data_1006 : _GEN_4077; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4079 = 10'h3ef == _dirty_T_1 ? cache_data_1007 : _GEN_4078; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4080 = 10'h3f0 == _dirty_T_1 ? cache_data_1008 : _GEN_4079; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4081 = 10'h3f1 == _dirty_T_1 ? cache_data_1009 : _GEN_4080; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4082 = 10'h3f2 == _dirty_T_1 ? cache_data_1010 : _GEN_4081; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4083 = 10'h3f3 == _dirty_T_1 ? cache_data_1011 : _GEN_4082; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4084 = 10'h3f4 == _dirty_T_1 ? cache_data_1012 : _GEN_4083; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4085 = 10'h3f5 == _dirty_T_1 ? cache_data_1013 : _GEN_4084; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4086 = 10'h3f6 == _dirty_T_1 ? cache_data_1014 : _GEN_4085; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4087 = 10'h3f7 == _dirty_T_1 ? cache_data_1015 : _GEN_4086; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4088 = 10'h3f8 == _dirty_T_1 ? cache_data_1016 : _GEN_4087; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4089 = 10'h3f9 == _dirty_T_1 ? cache_data_1017 : _GEN_4088; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4090 = 10'h3fa == _dirty_T_1 ? cache_data_1018 : _GEN_4089; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4091 = 10'h3fb == _dirty_T_1 ? cache_data_1019 : _GEN_4090; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4092 = 10'h3fc == _dirty_T_1 ? cache_data_1020 : _GEN_4091; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4093 = 10'h3fd == _dirty_T_1 ? cache_data_1021 : _GEN_4092; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4094 = 10'h3fe == _dirty_T_1 ? cache_data_1022 : _GEN_4093; // @[icache.scala 51:{42,42}]
  wire [184:0] _GEN_4095 = 10'h3ff == _dirty_T_1 ? cache_data_1023 : _GEN_4094; // @[icache.scala 51:{42,42}]
  wire  dirty = _GEN_4095[184:183] == 2'h3; // @[icache.scala 51:53]
  wire [1:0] _GEN_4097 = dirty ? 2'h2 : 2'h3; // @[icache.scala 65:27 66:17 68:17]
  wire [1:0] _GEN_4098 = hit ? 2'h1 : _GEN_4097; // @[icache.scala 63:19 64:17]
  wire [1:0] _GEN_4099 = io_valid ? _GEN_4098 : 2'h0; // @[icache.scala 62:22 71:15]
  wire [1:0] _GEN_4100 = io_rd_rdy ? 2'h3 : 2'h2; // @[icache.scala 75:23 76:15 78:15]
  wire [1:0] _GEN_4101 = io_inst_sram_data_ok ? 2'h1 : 2'h3; // @[icache.scala 82:34 83:15 85:15]
  wire [1:0] _GEN_4102 = 2'h3 == state ? _GEN_4101 : state; // @[icache.scala 53:17 23:67]
  wire [1:0] _GEN_4103 = 2'h2 == state ? _GEN_4100 : _GEN_4102; // @[icache.scala 53:17]
  wire  _T_5 = lookup & hit; // @[icache.scala 103:15]
  wire [184:0] _GEN_6158 = reset ? 185'h0 : cache_data_0; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6159 = reset ? 185'h0 : cache_data_1; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6160 = reset ? 185'h0 : cache_data_2; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6161 = reset ? 185'h0 : cache_data_3; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6162 = reset ? 185'h0 : cache_data_4; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6163 = reset ? 185'h0 : cache_data_5; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6164 = reset ? 185'h0 : cache_data_6; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6165 = reset ? 185'h0 : cache_data_7; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6166 = reset ? 185'h0 : cache_data_8; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6167 = reset ? 185'h0 : cache_data_9; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6168 = reset ? 185'h0 : cache_data_10; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6169 = reset ? 185'h0 : cache_data_11; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6170 = reset ? 185'h0 : cache_data_12; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6171 = reset ? 185'h0 : cache_data_13; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6172 = reset ? 185'h0 : cache_data_14; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6173 = reset ? 185'h0 : cache_data_15; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6174 = reset ? 185'h0 : cache_data_16; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6175 = reset ? 185'h0 : cache_data_17; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6176 = reset ? 185'h0 : cache_data_18; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6177 = reset ? 185'h0 : cache_data_19; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6178 = reset ? 185'h0 : cache_data_20; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6179 = reset ? 185'h0 : cache_data_21; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6180 = reset ? 185'h0 : cache_data_22; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6181 = reset ? 185'h0 : cache_data_23; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6182 = reset ? 185'h0 : cache_data_24; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6183 = reset ? 185'h0 : cache_data_25; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6184 = reset ? 185'h0 : cache_data_26; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6185 = reset ? 185'h0 : cache_data_27; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6186 = reset ? 185'h0 : cache_data_28; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6187 = reset ? 185'h0 : cache_data_29; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6188 = reset ? 185'h0 : cache_data_30; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6189 = reset ? 185'h0 : cache_data_31; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6190 = reset ? 185'h0 : cache_data_32; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6191 = reset ? 185'h0 : cache_data_33; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6192 = reset ? 185'h0 : cache_data_34; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6193 = reset ? 185'h0 : cache_data_35; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6194 = reset ? 185'h0 : cache_data_36; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6195 = reset ? 185'h0 : cache_data_37; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6196 = reset ? 185'h0 : cache_data_38; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6197 = reset ? 185'h0 : cache_data_39; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6198 = reset ? 185'h0 : cache_data_40; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6199 = reset ? 185'h0 : cache_data_41; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6200 = reset ? 185'h0 : cache_data_42; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6201 = reset ? 185'h0 : cache_data_43; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6202 = reset ? 185'h0 : cache_data_44; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6203 = reset ? 185'h0 : cache_data_45; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6204 = reset ? 185'h0 : cache_data_46; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6205 = reset ? 185'h0 : cache_data_47; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6206 = reset ? 185'h0 : cache_data_48; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6207 = reset ? 185'h0 : cache_data_49; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6208 = reset ? 185'h0 : cache_data_50; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6209 = reset ? 185'h0 : cache_data_51; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6210 = reset ? 185'h0 : cache_data_52; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6211 = reset ? 185'h0 : cache_data_53; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6212 = reset ? 185'h0 : cache_data_54; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6213 = reset ? 185'h0 : cache_data_55; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6214 = reset ? 185'h0 : cache_data_56; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6215 = reset ? 185'h0 : cache_data_57; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6216 = reset ? 185'h0 : cache_data_58; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6217 = reset ? 185'h0 : cache_data_59; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6218 = reset ? 185'h0 : cache_data_60; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6219 = reset ? 185'h0 : cache_data_61; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6220 = reset ? 185'h0 : cache_data_62; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6221 = reset ? 185'h0 : cache_data_63; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6222 = reset ? 185'h0 : cache_data_64; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6223 = reset ? 185'h0 : cache_data_65; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6224 = reset ? 185'h0 : cache_data_66; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6225 = reset ? 185'h0 : cache_data_67; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6226 = reset ? 185'h0 : cache_data_68; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6227 = reset ? 185'h0 : cache_data_69; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6228 = reset ? 185'h0 : cache_data_70; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6229 = reset ? 185'h0 : cache_data_71; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6230 = reset ? 185'h0 : cache_data_72; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6231 = reset ? 185'h0 : cache_data_73; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6232 = reset ? 185'h0 : cache_data_74; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6233 = reset ? 185'h0 : cache_data_75; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6234 = reset ? 185'h0 : cache_data_76; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6235 = reset ? 185'h0 : cache_data_77; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6236 = reset ? 185'h0 : cache_data_78; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6237 = reset ? 185'h0 : cache_data_79; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6238 = reset ? 185'h0 : cache_data_80; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6239 = reset ? 185'h0 : cache_data_81; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6240 = reset ? 185'h0 : cache_data_82; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6241 = reset ? 185'h0 : cache_data_83; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6242 = reset ? 185'h0 : cache_data_84; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6243 = reset ? 185'h0 : cache_data_85; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6244 = reset ? 185'h0 : cache_data_86; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6245 = reset ? 185'h0 : cache_data_87; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6246 = reset ? 185'h0 : cache_data_88; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6247 = reset ? 185'h0 : cache_data_89; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6248 = reset ? 185'h0 : cache_data_90; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6249 = reset ? 185'h0 : cache_data_91; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6250 = reset ? 185'h0 : cache_data_92; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6251 = reset ? 185'h0 : cache_data_93; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6252 = reset ? 185'h0 : cache_data_94; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6253 = reset ? 185'h0 : cache_data_95; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6254 = reset ? 185'h0 : cache_data_96; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6255 = reset ? 185'h0 : cache_data_97; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6256 = reset ? 185'h0 : cache_data_98; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6257 = reset ? 185'h0 : cache_data_99; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6258 = reset ? 185'h0 : cache_data_100; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6259 = reset ? 185'h0 : cache_data_101; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6260 = reset ? 185'h0 : cache_data_102; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6261 = reset ? 185'h0 : cache_data_103; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6262 = reset ? 185'h0 : cache_data_104; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6263 = reset ? 185'h0 : cache_data_105; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6264 = reset ? 185'h0 : cache_data_106; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6265 = reset ? 185'h0 : cache_data_107; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6266 = reset ? 185'h0 : cache_data_108; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6267 = reset ? 185'h0 : cache_data_109; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6268 = reset ? 185'h0 : cache_data_110; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6269 = reset ? 185'h0 : cache_data_111; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6270 = reset ? 185'h0 : cache_data_112; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6271 = reset ? 185'h0 : cache_data_113; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6272 = reset ? 185'h0 : cache_data_114; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6273 = reset ? 185'h0 : cache_data_115; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6274 = reset ? 185'h0 : cache_data_116; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6275 = reset ? 185'h0 : cache_data_117; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6276 = reset ? 185'h0 : cache_data_118; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6277 = reset ? 185'h0 : cache_data_119; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6278 = reset ? 185'h0 : cache_data_120; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6279 = reset ? 185'h0 : cache_data_121; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6280 = reset ? 185'h0 : cache_data_122; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6281 = reset ? 185'h0 : cache_data_123; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6282 = reset ? 185'h0 : cache_data_124; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6283 = reset ? 185'h0 : cache_data_125; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6284 = reset ? 185'h0 : cache_data_126; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6285 = reset ? 185'h0 : cache_data_127; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6286 = reset ? 185'h0 : cache_data_128; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6287 = reset ? 185'h0 : cache_data_129; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6288 = reset ? 185'h0 : cache_data_130; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6289 = reset ? 185'h0 : cache_data_131; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6290 = reset ? 185'h0 : cache_data_132; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6291 = reset ? 185'h0 : cache_data_133; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6292 = reset ? 185'h0 : cache_data_134; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6293 = reset ? 185'h0 : cache_data_135; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6294 = reset ? 185'h0 : cache_data_136; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6295 = reset ? 185'h0 : cache_data_137; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6296 = reset ? 185'h0 : cache_data_138; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6297 = reset ? 185'h0 : cache_data_139; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6298 = reset ? 185'h0 : cache_data_140; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6299 = reset ? 185'h0 : cache_data_141; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6300 = reset ? 185'h0 : cache_data_142; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6301 = reset ? 185'h0 : cache_data_143; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6302 = reset ? 185'h0 : cache_data_144; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6303 = reset ? 185'h0 : cache_data_145; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6304 = reset ? 185'h0 : cache_data_146; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6305 = reset ? 185'h0 : cache_data_147; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6306 = reset ? 185'h0 : cache_data_148; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6307 = reset ? 185'h0 : cache_data_149; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6308 = reset ? 185'h0 : cache_data_150; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6309 = reset ? 185'h0 : cache_data_151; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6310 = reset ? 185'h0 : cache_data_152; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6311 = reset ? 185'h0 : cache_data_153; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6312 = reset ? 185'h0 : cache_data_154; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6313 = reset ? 185'h0 : cache_data_155; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6314 = reset ? 185'h0 : cache_data_156; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6315 = reset ? 185'h0 : cache_data_157; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6316 = reset ? 185'h0 : cache_data_158; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6317 = reset ? 185'h0 : cache_data_159; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6318 = reset ? 185'h0 : cache_data_160; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6319 = reset ? 185'h0 : cache_data_161; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6320 = reset ? 185'h0 : cache_data_162; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6321 = reset ? 185'h0 : cache_data_163; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6322 = reset ? 185'h0 : cache_data_164; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6323 = reset ? 185'h0 : cache_data_165; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6324 = reset ? 185'h0 : cache_data_166; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6325 = reset ? 185'h0 : cache_data_167; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6326 = reset ? 185'h0 : cache_data_168; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6327 = reset ? 185'h0 : cache_data_169; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6328 = reset ? 185'h0 : cache_data_170; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6329 = reset ? 185'h0 : cache_data_171; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6330 = reset ? 185'h0 : cache_data_172; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6331 = reset ? 185'h0 : cache_data_173; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6332 = reset ? 185'h0 : cache_data_174; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6333 = reset ? 185'h0 : cache_data_175; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6334 = reset ? 185'h0 : cache_data_176; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6335 = reset ? 185'h0 : cache_data_177; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6336 = reset ? 185'h0 : cache_data_178; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6337 = reset ? 185'h0 : cache_data_179; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6338 = reset ? 185'h0 : cache_data_180; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6339 = reset ? 185'h0 : cache_data_181; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6340 = reset ? 185'h0 : cache_data_182; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6341 = reset ? 185'h0 : cache_data_183; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6342 = reset ? 185'h0 : cache_data_184; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6343 = reset ? 185'h0 : cache_data_185; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6344 = reset ? 185'h0 : cache_data_186; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6345 = reset ? 185'h0 : cache_data_187; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6346 = reset ? 185'h0 : cache_data_188; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6347 = reset ? 185'h0 : cache_data_189; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6348 = reset ? 185'h0 : cache_data_190; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6349 = reset ? 185'h0 : cache_data_191; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6350 = reset ? 185'h0 : cache_data_192; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6351 = reset ? 185'h0 : cache_data_193; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6352 = reset ? 185'h0 : cache_data_194; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6353 = reset ? 185'h0 : cache_data_195; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6354 = reset ? 185'h0 : cache_data_196; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6355 = reset ? 185'h0 : cache_data_197; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6356 = reset ? 185'h0 : cache_data_198; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6357 = reset ? 185'h0 : cache_data_199; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6358 = reset ? 185'h0 : cache_data_200; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6359 = reset ? 185'h0 : cache_data_201; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6360 = reset ? 185'h0 : cache_data_202; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6361 = reset ? 185'h0 : cache_data_203; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6362 = reset ? 185'h0 : cache_data_204; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6363 = reset ? 185'h0 : cache_data_205; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6364 = reset ? 185'h0 : cache_data_206; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6365 = reset ? 185'h0 : cache_data_207; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6366 = reset ? 185'h0 : cache_data_208; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6367 = reset ? 185'h0 : cache_data_209; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6368 = reset ? 185'h0 : cache_data_210; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6369 = reset ? 185'h0 : cache_data_211; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6370 = reset ? 185'h0 : cache_data_212; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6371 = reset ? 185'h0 : cache_data_213; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6372 = reset ? 185'h0 : cache_data_214; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6373 = reset ? 185'h0 : cache_data_215; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6374 = reset ? 185'h0 : cache_data_216; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6375 = reset ? 185'h0 : cache_data_217; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6376 = reset ? 185'h0 : cache_data_218; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6377 = reset ? 185'h0 : cache_data_219; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6378 = reset ? 185'h0 : cache_data_220; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6379 = reset ? 185'h0 : cache_data_221; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6380 = reset ? 185'h0 : cache_data_222; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6381 = reset ? 185'h0 : cache_data_223; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6382 = reset ? 185'h0 : cache_data_224; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6383 = reset ? 185'h0 : cache_data_225; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6384 = reset ? 185'h0 : cache_data_226; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6385 = reset ? 185'h0 : cache_data_227; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6386 = reset ? 185'h0 : cache_data_228; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6387 = reset ? 185'h0 : cache_data_229; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6388 = reset ? 185'h0 : cache_data_230; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6389 = reset ? 185'h0 : cache_data_231; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6390 = reset ? 185'h0 : cache_data_232; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6391 = reset ? 185'h0 : cache_data_233; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6392 = reset ? 185'h0 : cache_data_234; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6393 = reset ? 185'h0 : cache_data_235; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6394 = reset ? 185'h0 : cache_data_236; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6395 = reset ? 185'h0 : cache_data_237; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6396 = reset ? 185'h0 : cache_data_238; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6397 = reset ? 185'h0 : cache_data_239; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6398 = reset ? 185'h0 : cache_data_240; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6399 = reset ? 185'h0 : cache_data_241; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6400 = reset ? 185'h0 : cache_data_242; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6401 = reset ? 185'h0 : cache_data_243; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6402 = reset ? 185'h0 : cache_data_244; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6403 = reset ? 185'h0 : cache_data_245; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6404 = reset ? 185'h0 : cache_data_246; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6405 = reset ? 185'h0 : cache_data_247; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6406 = reset ? 185'h0 : cache_data_248; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6407 = reset ? 185'h0 : cache_data_249; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6408 = reset ? 185'h0 : cache_data_250; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6409 = reset ? 185'h0 : cache_data_251; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6410 = reset ? 185'h0 : cache_data_252; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6411 = reset ? 185'h0 : cache_data_253; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6412 = reset ? 185'h0 : cache_data_254; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6413 = reset ? 185'h0 : cache_data_255; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6414 = reset ? 185'h0 : cache_data_256; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6415 = reset ? 185'h0 : cache_data_257; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6416 = reset ? 185'h0 : cache_data_258; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6417 = reset ? 185'h0 : cache_data_259; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6418 = reset ? 185'h0 : cache_data_260; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6419 = reset ? 185'h0 : cache_data_261; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6420 = reset ? 185'h0 : cache_data_262; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6421 = reset ? 185'h0 : cache_data_263; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6422 = reset ? 185'h0 : cache_data_264; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6423 = reset ? 185'h0 : cache_data_265; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6424 = reset ? 185'h0 : cache_data_266; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6425 = reset ? 185'h0 : cache_data_267; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6426 = reset ? 185'h0 : cache_data_268; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6427 = reset ? 185'h0 : cache_data_269; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6428 = reset ? 185'h0 : cache_data_270; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6429 = reset ? 185'h0 : cache_data_271; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6430 = reset ? 185'h0 : cache_data_272; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6431 = reset ? 185'h0 : cache_data_273; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6432 = reset ? 185'h0 : cache_data_274; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6433 = reset ? 185'h0 : cache_data_275; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6434 = reset ? 185'h0 : cache_data_276; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6435 = reset ? 185'h0 : cache_data_277; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6436 = reset ? 185'h0 : cache_data_278; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6437 = reset ? 185'h0 : cache_data_279; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6438 = reset ? 185'h0 : cache_data_280; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6439 = reset ? 185'h0 : cache_data_281; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6440 = reset ? 185'h0 : cache_data_282; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6441 = reset ? 185'h0 : cache_data_283; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6442 = reset ? 185'h0 : cache_data_284; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6443 = reset ? 185'h0 : cache_data_285; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6444 = reset ? 185'h0 : cache_data_286; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6445 = reset ? 185'h0 : cache_data_287; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6446 = reset ? 185'h0 : cache_data_288; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6447 = reset ? 185'h0 : cache_data_289; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6448 = reset ? 185'h0 : cache_data_290; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6449 = reset ? 185'h0 : cache_data_291; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6450 = reset ? 185'h0 : cache_data_292; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6451 = reset ? 185'h0 : cache_data_293; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6452 = reset ? 185'h0 : cache_data_294; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6453 = reset ? 185'h0 : cache_data_295; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6454 = reset ? 185'h0 : cache_data_296; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6455 = reset ? 185'h0 : cache_data_297; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6456 = reset ? 185'h0 : cache_data_298; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6457 = reset ? 185'h0 : cache_data_299; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6458 = reset ? 185'h0 : cache_data_300; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6459 = reset ? 185'h0 : cache_data_301; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6460 = reset ? 185'h0 : cache_data_302; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6461 = reset ? 185'h0 : cache_data_303; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6462 = reset ? 185'h0 : cache_data_304; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6463 = reset ? 185'h0 : cache_data_305; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6464 = reset ? 185'h0 : cache_data_306; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6465 = reset ? 185'h0 : cache_data_307; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6466 = reset ? 185'h0 : cache_data_308; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6467 = reset ? 185'h0 : cache_data_309; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6468 = reset ? 185'h0 : cache_data_310; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6469 = reset ? 185'h0 : cache_data_311; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6470 = reset ? 185'h0 : cache_data_312; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6471 = reset ? 185'h0 : cache_data_313; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6472 = reset ? 185'h0 : cache_data_314; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6473 = reset ? 185'h0 : cache_data_315; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6474 = reset ? 185'h0 : cache_data_316; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6475 = reset ? 185'h0 : cache_data_317; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6476 = reset ? 185'h0 : cache_data_318; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6477 = reset ? 185'h0 : cache_data_319; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6478 = reset ? 185'h0 : cache_data_320; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6479 = reset ? 185'h0 : cache_data_321; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6480 = reset ? 185'h0 : cache_data_322; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6481 = reset ? 185'h0 : cache_data_323; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6482 = reset ? 185'h0 : cache_data_324; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6483 = reset ? 185'h0 : cache_data_325; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6484 = reset ? 185'h0 : cache_data_326; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6485 = reset ? 185'h0 : cache_data_327; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6486 = reset ? 185'h0 : cache_data_328; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6487 = reset ? 185'h0 : cache_data_329; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6488 = reset ? 185'h0 : cache_data_330; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6489 = reset ? 185'h0 : cache_data_331; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6490 = reset ? 185'h0 : cache_data_332; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6491 = reset ? 185'h0 : cache_data_333; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6492 = reset ? 185'h0 : cache_data_334; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6493 = reset ? 185'h0 : cache_data_335; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6494 = reset ? 185'h0 : cache_data_336; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6495 = reset ? 185'h0 : cache_data_337; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6496 = reset ? 185'h0 : cache_data_338; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6497 = reset ? 185'h0 : cache_data_339; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6498 = reset ? 185'h0 : cache_data_340; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6499 = reset ? 185'h0 : cache_data_341; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6500 = reset ? 185'h0 : cache_data_342; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6501 = reset ? 185'h0 : cache_data_343; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6502 = reset ? 185'h0 : cache_data_344; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6503 = reset ? 185'h0 : cache_data_345; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6504 = reset ? 185'h0 : cache_data_346; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6505 = reset ? 185'h0 : cache_data_347; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6506 = reset ? 185'h0 : cache_data_348; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6507 = reset ? 185'h0 : cache_data_349; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6508 = reset ? 185'h0 : cache_data_350; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6509 = reset ? 185'h0 : cache_data_351; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6510 = reset ? 185'h0 : cache_data_352; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6511 = reset ? 185'h0 : cache_data_353; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6512 = reset ? 185'h0 : cache_data_354; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6513 = reset ? 185'h0 : cache_data_355; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6514 = reset ? 185'h0 : cache_data_356; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6515 = reset ? 185'h0 : cache_data_357; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6516 = reset ? 185'h0 : cache_data_358; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6517 = reset ? 185'h0 : cache_data_359; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6518 = reset ? 185'h0 : cache_data_360; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6519 = reset ? 185'h0 : cache_data_361; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6520 = reset ? 185'h0 : cache_data_362; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6521 = reset ? 185'h0 : cache_data_363; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6522 = reset ? 185'h0 : cache_data_364; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6523 = reset ? 185'h0 : cache_data_365; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6524 = reset ? 185'h0 : cache_data_366; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6525 = reset ? 185'h0 : cache_data_367; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6526 = reset ? 185'h0 : cache_data_368; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6527 = reset ? 185'h0 : cache_data_369; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6528 = reset ? 185'h0 : cache_data_370; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6529 = reset ? 185'h0 : cache_data_371; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6530 = reset ? 185'h0 : cache_data_372; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6531 = reset ? 185'h0 : cache_data_373; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6532 = reset ? 185'h0 : cache_data_374; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6533 = reset ? 185'h0 : cache_data_375; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6534 = reset ? 185'h0 : cache_data_376; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6535 = reset ? 185'h0 : cache_data_377; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6536 = reset ? 185'h0 : cache_data_378; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6537 = reset ? 185'h0 : cache_data_379; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6538 = reset ? 185'h0 : cache_data_380; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6539 = reset ? 185'h0 : cache_data_381; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6540 = reset ? 185'h0 : cache_data_382; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6541 = reset ? 185'h0 : cache_data_383; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6542 = reset ? 185'h0 : cache_data_384; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6543 = reset ? 185'h0 : cache_data_385; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6544 = reset ? 185'h0 : cache_data_386; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6545 = reset ? 185'h0 : cache_data_387; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6546 = reset ? 185'h0 : cache_data_388; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6547 = reset ? 185'h0 : cache_data_389; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6548 = reset ? 185'h0 : cache_data_390; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6549 = reset ? 185'h0 : cache_data_391; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6550 = reset ? 185'h0 : cache_data_392; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6551 = reset ? 185'h0 : cache_data_393; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6552 = reset ? 185'h0 : cache_data_394; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6553 = reset ? 185'h0 : cache_data_395; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6554 = reset ? 185'h0 : cache_data_396; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6555 = reset ? 185'h0 : cache_data_397; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6556 = reset ? 185'h0 : cache_data_398; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6557 = reset ? 185'h0 : cache_data_399; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6558 = reset ? 185'h0 : cache_data_400; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6559 = reset ? 185'h0 : cache_data_401; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6560 = reset ? 185'h0 : cache_data_402; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6561 = reset ? 185'h0 : cache_data_403; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6562 = reset ? 185'h0 : cache_data_404; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6563 = reset ? 185'h0 : cache_data_405; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6564 = reset ? 185'h0 : cache_data_406; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6565 = reset ? 185'h0 : cache_data_407; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6566 = reset ? 185'h0 : cache_data_408; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6567 = reset ? 185'h0 : cache_data_409; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6568 = reset ? 185'h0 : cache_data_410; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6569 = reset ? 185'h0 : cache_data_411; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6570 = reset ? 185'h0 : cache_data_412; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6571 = reset ? 185'h0 : cache_data_413; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6572 = reset ? 185'h0 : cache_data_414; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6573 = reset ? 185'h0 : cache_data_415; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6574 = reset ? 185'h0 : cache_data_416; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6575 = reset ? 185'h0 : cache_data_417; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6576 = reset ? 185'h0 : cache_data_418; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6577 = reset ? 185'h0 : cache_data_419; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6578 = reset ? 185'h0 : cache_data_420; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6579 = reset ? 185'h0 : cache_data_421; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6580 = reset ? 185'h0 : cache_data_422; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6581 = reset ? 185'h0 : cache_data_423; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6582 = reset ? 185'h0 : cache_data_424; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6583 = reset ? 185'h0 : cache_data_425; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6584 = reset ? 185'h0 : cache_data_426; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6585 = reset ? 185'h0 : cache_data_427; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6586 = reset ? 185'h0 : cache_data_428; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6587 = reset ? 185'h0 : cache_data_429; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6588 = reset ? 185'h0 : cache_data_430; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6589 = reset ? 185'h0 : cache_data_431; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6590 = reset ? 185'h0 : cache_data_432; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6591 = reset ? 185'h0 : cache_data_433; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6592 = reset ? 185'h0 : cache_data_434; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6593 = reset ? 185'h0 : cache_data_435; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6594 = reset ? 185'h0 : cache_data_436; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6595 = reset ? 185'h0 : cache_data_437; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6596 = reset ? 185'h0 : cache_data_438; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6597 = reset ? 185'h0 : cache_data_439; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6598 = reset ? 185'h0 : cache_data_440; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6599 = reset ? 185'h0 : cache_data_441; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6600 = reset ? 185'h0 : cache_data_442; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6601 = reset ? 185'h0 : cache_data_443; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6602 = reset ? 185'h0 : cache_data_444; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6603 = reset ? 185'h0 : cache_data_445; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6604 = reset ? 185'h0 : cache_data_446; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6605 = reset ? 185'h0 : cache_data_447; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6606 = reset ? 185'h0 : cache_data_448; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6607 = reset ? 185'h0 : cache_data_449; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6608 = reset ? 185'h0 : cache_data_450; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6609 = reset ? 185'h0 : cache_data_451; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6610 = reset ? 185'h0 : cache_data_452; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6611 = reset ? 185'h0 : cache_data_453; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6612 = reset ? 185'h0 : cache_data_454; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6613 = reset ? 185'h0 : cache_data_455; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6614 = reset ? 185'h0 : cache_data_456; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6615 = reset ? 185'h0 : cache_data_457; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6616 = reset ? 185'h0 : cache_data_458; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6617 = reset ? 185'h0 : cache_data_459; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6618 = reset ? 185'h0 : cache_data_460; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6619 = reset ? 185'h0 : cache_data_461; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6620 = reset ? 185'h0 : cache_data_462; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6621 = reset ? 185'h0 : cache_data_463; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6622 = reset ? 185'h0 : cache_data_464; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6623 = reset ? 185'h0 : cache_data_465; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6624 = reset ? 185'h0 : cache_data_466; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6625 = reset ? 185'h0 : cache_data_467; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6626 = reset ? 185'h0 : cache_data_468; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6627 = reset ? 185'h0 : cache_data_469; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6628 = reset ? 185'h0 : cache_data_470; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6629 = reset ? 185'h0 : cache_data_471; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6630 = reset ? 185'h0 : cache_data_472; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6631 = reset ? 185'h0 : cache_data_473; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6632 = reset ? 185'h0 : cache_data_474; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6633 = reset ? 185'h0 : cache_data_475; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6634 = reset ? 185'h0 : cache_data_476; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6635 = reset ? 185'h0 : cache_data_477; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6636 = reset ? 185'h0 : cache_data_478; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6637 = reset ? 185'h0 : cache_data_479; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6638 = reset ? 185'h0 : cache_data_480; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6639 = reset ? 185'h0 : cache_data_481; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6640 = reset ? 185'h0 : cache_data_482; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6641 = reset ? 185'h0 : cache_data_483; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6642 = reset ? 185'h0 : cache_data_484; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6643 = reset ? 185'h0 : cache_data_485; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6644 = reset ? 185'h0 : cache_data_486; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6645 = reset ? 185'h0 : cache_data_487; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6646 = reset ? 185'h0 : cache_data_488; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6647 = reset ? 185'h0 : cache_data_489; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6648 = reset ? 185'h0 : cache_data_490; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6649 = reset ? 185'h0 : cache_data_491; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6650 = reset ? 185'h0 : cache_data_492; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6651 = reset ? 185'h0 : cache_data_493; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6652 = reset ? 185'h0 : cache_data_494; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6653 = reset ? 185'h0 : cache_data_495; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6654 = reset ? 185'h0 : cache_data_496; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6655 = reset ? 185'h0 : cache_data_497; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6656 = reset ? 185'h0 : cache_data_498; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6657 = reset ? 185'h0 : cache_data_499; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6658 = reset ? 185'h0 : cache_data_500; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6659 = reset ? 185'h0 : cache_data_501; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6660 = reset ? 185'h0 : cache_data_502; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6661 = reset ? 185'h0 : cache_data_503; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6662 = reset ? 185'h0 : cache_data_504; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6663 = reset ? 185'h0 : cache_data_505; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6664 = reset ? 185'h0 : cache_data_506; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6665 = reset ? 185'h0 : cache_data_507; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6666 = reset ? 185'h0 : cache_data_508; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6667 = reset ? 185'h0 : cache_data_509; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6668 = reset ? 185'h0 : cache_data_510; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6669 = reset ? 185'h0 : cache_data_511; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6670 = reset ? 185'h0 : cache_data_512; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6671 = reset ? 185'h0 : cache_data_513; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6672 = reset ? 185'h0 : cache_data_514; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6673 = reset ? 185'h0 : cache_data_515; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6674 = reset ? 185'h0 : cache_data_516; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6675 = reset ? 185'h0 : cache_data_517; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6676 = reset ? 185'h0 : cache_data_518; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6677 = reset ? 185'h0 : cache_data_519; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6678 = reset ? 185'h0 : cache_data_520; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6679 = reset ? 185'h0 : cache_data_521; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6680 = reset ? 185'h0 : cache_data_522; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6681 = reset ? 185'h0 : cache_data_523; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6682 = reset ? 185'h0 : cache_data_524; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6683 = reset ? 185'h0 : cache_data_525; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6684 = reset ? 185'h0 : cache_data_526; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6685 = reset ? 185'h0 : cache_data_527; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6686 = reset ? 185'h0 : cache_data_528; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6687 = reset ? 185'h0 : cache_data_529; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6688 = reset ? 185'h0 : cache_data_530; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6689 = reset ? 185'h0 : cache_data_531; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6690 = reset ? 185'h0 : cache_data_532; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6691 = reset ? 185'h0 : cache_data_533; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6692 = reset ? 185'h0 : cache_data_534; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6693 = reset ? 185'h0 : cache_data_535; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6694 = reset ? 185'h0 : cache_data_536; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6695 = reset ? 185'h0 : cache_data_537; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6696 = reset ? 185'h0 : cache_data_538; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6697 = reset ? 185'h0 : cache_data_539; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6698 = reset ? 185'h0 : cache_data_540; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6699 = reset ? 185'h0 : cache_data_541; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6700 = reset ? 185'h0 : cache_data_542; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6701 = reset ? 185'h0 : cache_data_543; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6702 = reset ? 185'h0 : cache_data_544; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6703 = reset ? 185'h0 : cache_data_545; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6704 = reset ? 185'h0 : cache_data_546; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6705 = reset ? 185'h0 : cache_data_547; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6706 = reset ? 185'h0 : cache_data_548; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6707 = reset ? 185'h0 : cache_data_549; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6708 = reset ? 185'h0 : cache_data_550; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6709 = reset ? 185'h0 : cache_data_551; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6710 = reset ? 185'h0 : cache_data_552; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6711 = reset ? 185'h0 : cache_data_553; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6712 = reset ? 185'h0 : cache_data_554; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6713 = reset ? 185'h0 : cache_data_555; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6714 = reset ? 185'h0 : cache_data_556; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6715 = reset ? 185'h0 : cache_data_557; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6716 = reset ? 185'h0 : cache_data_558; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6717 = reset ? 185'h0 : cache_data_559; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6718 = reset ? 185'h0 : cache_data_560; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6719 = reset ? 185'h0 : cache_data_561; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6720 = reset ? 185'h0 : cache_data_562; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6721 = reset ? 185'h0 : cache_data_563; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6722 = reset ? 185'h0 : cache_data_564; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6723 = reset ? 185'h0 : cache_data_565; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6724 = reset ? 185'h0 : cache_data_566; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6725 = reset ? 185'h0 : cache_data_567; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6726 = reset ? 185'h0 : cache_data_568; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6727 = reset ? 185'h0 : cache_data_569; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6728 = reset ? 185'h0 : cache_data_570; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6729 = reset ? 185'h0 : cache_data_571; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6730 = reset ? 185'h0 : cache_data_572; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6731 = reset ? 185'h0 : cache_data_573; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6732 = reset ? 185'h0 : cache_data_574; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6733 = reset ? 185'h0 : cache_data_575; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6734 = reset ? 185'h0 : cache_data_576; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6735 = reset ? 185'h0 : cache_data_577; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6736 = reset ? 185'h0 : cache_data_578; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6737 = reset ? 185'h0 : cache_data_579; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6738 = reset ? 185'h0 : cache_data_580; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6739 = reset ? 185'h0 : cache_data_581; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6740 = reset ? 185'h0 : cache_data_582; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6741 = reset ? 185'h0 : cache_data_583; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6742 = reset ? 185'h0 : cache_data_584; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6743 = reset ? 185'h0 : cache_data_585; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6744 = reset ? 185'h0 : cache_data_586; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6745 = reset ? 185'h0 : cache_data_587; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6746 = reset ? 185'h0 : cache_data_588; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6747 = reset ? 185'h0 : cache_data_589; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6748 = reset ? 185'h0 : cache_data_590; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6749 = reset ? 185'h0 : cache_data_591; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6750 = reset ? 185'h0 : cache_data_592; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6751 = reset ? 185'h0 : cache_data_593; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6752 = reset ? 185'h0 : cache_data_594; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6753 = reset ? 185'h0 : cache_data_595; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6754 = reset ? 185'h0 : cache_data_596; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6755 = reset ? 185'h0 : cache_data_597; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6756 = reset ? 185'h0 : cache_data_598; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6757 = reset ? 185'h0 : cache_data_599; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6758 = reset ? 185'h0 : cache_data_600; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6759 = reset ? 185'h0 : cache_data_601; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6760 = reset ? 185'h0 : cache_data_602; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6761 = reset ? 185'h0 : cache_data_603; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6762 = reset ? 185'h0 : cache_data_604; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6763 = reset ? 185'h0 : cache_data_605; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6764 = reset ? 185'h0 : cache_data_606; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6765 = reset ? 185'h0 : cache_data_607; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6766 = reset ? 185'h0 : cache_data_608; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6767 = reset ? 185'h0 : cache_data_609; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6768 = reset ? 185'h0 : cache_data_610; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6769 = reset ? 185'h0 : cache_data_611; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6770 = reset ? 185'h0 : cache_data_612; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6771 = reset ? 185'h0 : cache_data_613; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6772 = reset ? 185'h0 : cache_data_614; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6773 = reset ? 185'h0 : cache_data_615; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6774 = reset ? 185'h0 : cache_data_616; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6775 = reset ? 185'h0 : cache_data_617; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6776 = reset ? 185'h0 : cache_data_618; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6777 = reset ? 185'h0 : cache_data_619; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6778 = reset ? 185'h0 : cache_data_620; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6779 = reset ? 185'h0 : cache_data_621; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6780 = reset ? 185'h0 : cache_data_622; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6781 = reset ? 185'h0 : cache_data_623; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6782 = reset ? 185'h0 : cache_data_624; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6783 = reset ? 185'h0 : cache_data_625; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6784 = reset ? 185'h0 : cache_data_626; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6785 = reset ? 185'h0 : cache_data_627; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6786 = reset ? 185'h0 : cache_data_628; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6787 = reset ? 185'h0 : cache_data_629; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6788 = reset ? 185'h0 : cache_data_630; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6789 = reset ? 185'h0 : cache_data_631; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6790 = reset ? 185'h0 : cache_data_632; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6791 = reset ? 185'h0 : cache_data_633; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6792 = reset ? 185'h0 : cache_data_634; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6793 = reset ? 185'h0 : cache_data_635; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6794 = reset ? 185'h0 : cache_data_636; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6795 = reset ? 185'h0 : cache_data_637; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6796 = reset ? 185'h0 : cache_data_638; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6797 = reset ? 185'h0 : cache_data_639; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6798 = reset ? 185'h0 : cache_data_640; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6799 = reset ? 185'h0 : cache_data_641; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6800 = reset ? 185'h0 : cache_data_642; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6801 = reset ? 185'h0 : cache_data_643; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6802 = reset ? 185'h0 : cache_data_644; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6803 = reset ? 185'h0 : cache_data_645; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6804 = reset ? 185'h0 : cache_data_646; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6805 = reset ? 185'h0 : cache_data_647; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6806 = reset ? 185'h0 : cache_data_648; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6807 = reset ? 185'h0 : cache_data_649; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6808 = reset ? 185'h0 : cache_data_650; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6809 = reset ? 185'h0 : cache_data_651; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6810 = reset ? 185'h0 : cache_data_652; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6811 = reset ? 185'h0 : cache_data_653; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6812 = reset ? 185'h0 : cache_data_654; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6813 = reset ? 185'h0 : cache_data_655; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6814 = reset ? 185'h0 : cache_data_656; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6815 = reset ? 185'h0 : cache_data_657; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6816 = reset ? 185'h0 : cache_data_658; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6817 = reset ? 185'h0 : cache_data_659; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6818 = reset ? 185'h0 : cache_data_660; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6819 = reset ? 185'h0 : cache_data_661; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6820 = reset ? 185'h0 : cache_data_662; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6821 = reset ? 185'h0 : cache_data_663; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6822 = reset ? 185'h0 : cache_data_664; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6823 = reset ? 185'h0 : cache_data_665; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6824 = reset ? 185'h0 : cache_data_666; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6825 = reset ? 185'h0 : cache_data_667; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6826 = reset ? 185'h0 : cache_data_668; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6827 = reset ? 185'h0 : cache_data_669; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6828 = reset ? 185'h0 : cache_data_670; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6829 = reset ? 185'h0 : cache_data_671; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6830 = reset ? 185'h0 : cache_data_672; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6831 = reset ? 185'h0 : cache_data_673; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6832 = reset ? 185'h0 : cache_data_674; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6833 = reset ? 185'h0 : cache_data_675; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6834 = reset ? 185'h0 : cache_data_676; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6835 = reset ? 185'h0 : cache_data_677; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6836 = reset ? 185'h0 : cache_data_678; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6837 = reset ? 185'h0 : cache_data_679; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6838 = reset ? 185'h0 : cache_data_680; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6839 = reset ? 185'h0 : cache_data_681; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6840 = reset ? 185'h0 : cache_data_682; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6841 = reset ? 185'h0 : cache_data_683; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6842 = reset ? 185'h0 : cache_data_684; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6843 = reset ? 185'h0 : cache_data_685; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6844 = reset ? 185'h0 : cache_data_686; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6845 = reset ? 185'h0 : cache_data_687; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6846 = reset ? 185'h0 : cache_data_688; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6847 = reset ? 185'h0 : cache_data_689; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6848 = reset ? 185'h0 : cache_data_690; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6849 = reset ? 185'h0 : cache_data_691; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6850 = reset ? 185'h0 : cache_data_692; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6851 = reset ? 185'h0 : cache_data_693; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6852 = reset ? 185'h0 : cache_data_694; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6853 = reset ? 185'h0 : cache_data_695; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6854 = reset ? 185'h0 : cache_data_696; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6855 = reset ? 185'h0 : cache_data_697; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6856 = reset ? 185'h0 : cache_data_698; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6857 = reset ? 185'h0 : cache_data_699; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6858 = reset ? 185'h0 : cache_data_700; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6859 = reset ? 185'h0 : cache_data_701; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6860 = reset ? 185'h0 : cache_data_702; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6861 = reset ? 185'h0 : cache_data_703; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6862 = reset ? 185'h0 : cache_data_704; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6863 = reset ? 185'h0 : cache_data_705; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6864 = reset ? 185'h0 : cache_data_706; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6865 = reset ? 185'h0 : cache_data_707; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6866 = reset ? 185'h0 : cache_data_708; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6867 = reset ? 185'h0 : cache_data_709; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6868 = reset ? 185'h0 : cache_data_710; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6869 = reset ? 185'h0 : cache_data_711; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6870 = reset ? 185'h0 : cache_data_712; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6871 = reset ? 185'h0 : cache_data_713; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6872 = reset ? 185'h0 : cache_data_714; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6873 = reset ? 185'h0 : cache_data_715; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6874 = reset ? 185'h0 : cache_data_716; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6875 = reset ? 185'h0 : cache_data_717; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6876 = reset ? 185'h0 : cache_data_718; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6877 = reset ? 185'h0 : cache_data_719; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6878 = reset ? 185'h0 : cache_data_720; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6879 = reset ? 185'h0 : cache_data_721; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6880 = reset ? 185'h0 : cache_data_722; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6881 = reset ? 185'h0 : cache_data_723; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6882 = reset ? 185'h0 : cache_data_724; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6883 = reset ? 185'h0 : cache_data_725; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6884 = reset ? 185'h0 : cache_data_726; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6885 = reset ? 185'h0 : cache_data_727; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6886 = reset ? 185'h0 : cache_data_728; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6887 = reset ? 185'h0 : cache_data_729; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6888 = reset ? 185'h0 : cache_data_730; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6889 = reset ? 185'h0 : cache_data_731; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6890 = reset ? 185'h0 : cache_data_732; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6891 = reset ? 185'h0 : cache_data_733; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6892 = reset ? 185'h0 : cache_data_734; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6893 = reset ? 185'h0 : cache_data_735; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6894 = reset ? 185'h0 : cache_data_736; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6895 = reset ? 185'h0 : cache_data_737; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6896 = reset ? 185'h0 : cache_data_738; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6897 = reset ? 185'h0 : cache_data_739; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6898 = reset ? 185'h0 : cache_data_740; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6899 = reset ? 185'h0 : cache_data_741; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6900 = reset ? 185'h0 : cache_data_742; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6901 = reset ? 185'h0 : cache_data_743; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6902 = reset ? 185'h0 : cache_data_744; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6903 = reset ? 185'h0 : cache_data_745; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6904 = reset ? 185'h0 : cache_data_746; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6905 = reset ? 185'h0 : cache_data_747; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6906 = reset ? 185'h0 : cache_data_748; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6907 = reset ? 185'h0 : cache_data_749; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6908 = reset ? 185'h0 : cache_data_750; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6909 = reset ? 185'h0 : cache_data_751; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6910 = reset ? 185'h0 : cache_data_752; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6911 = reset ? 185'h0 : cache_data_753; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6912 = reset ? 185'h0 : cache_data_754; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6913 = reset ? 185'h0 : cache_data_755; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6914 = reset ? 185'h0 : cache_data_756; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6915 = reset ? 185'h0 : cache_data_757; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6916 = reset ? 185'h0 : cache_data_758; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6917 = reset ? 185'h0 : cache_data_759; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6918 = reset ? 185'h0 : cache_data_760; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6919 = reset ? 185'h0 : cache_data_761; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6920 = reset ? 185'h0 : cache_data_762; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6921 = reset ? 185'h0 : cache_data_763; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6922 = reset ? 185'h0 : cache_data_764; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6923 = reset ? 185'h0 : cache_data_765; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6924 = reset ? 185'h0 : cache_data_766; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6925 = reset ? 185'h0 : cache_data_767; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6926 = reset ? 185'h0 : cache_data_768; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6927 = reset ? 185'h0 : cache_data_769; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6928 = reset ? 185'h0 : cache_data_770; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6929 = reset ? 185'h0 : cache_data_771; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6930 = reset ? 185'h0 : cache_data_772; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6931 = reset ? 185'h0 : cache_data_773; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6932 = reset ? 185'h0 : cache_data_774; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6933 = reset ? 185'h0 : cache_data_775; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6934 = reset ? 185'h0 : cache_data_776; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6935 = reset ? 185'h0 : cache_data_777; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6936 = reset ? 185'h0 : cache_data_778; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6937 = reset ? 185'h0 : cache_data_779; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6938 = reset ? 185'h0 : cache_data_780; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6939 = reset ? 185'h0 : cache_data_781; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6940 = reset ? 185'h0 : cache_data_782; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6941 = reset ? 185'h0 : cache_data_783; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6942 = reset ? 185'h0 : cache_data_784; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6943 = reset ? 185'h0 : cache_data_785; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6944 = reset ? 185'h0 : cache_data_786; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6945 = reset ? 185'h0 : cache_data_787; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6946 = reset ? 185'h0 : cache_data_788; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6947 = reset ? 185'h0 : cache_data_789; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6948 = reset ? 185'h0 : cache_data_790; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6949 = reset ? 185'h0 : cache_data_791; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6950 = reset ? 185'h0 : cache_data_792; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6951 = reset ? 185'h0 : cache_data_793; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6952 = reset ? 185'h0 : cache_data_794; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6953 = reset ? 185'h0 : cache_data_795; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6954 = reset ? 185'h0 : cache_data_796; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6955 = reset ? 185'h0 : cache_data_797; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6956 = reset ? 185'h0 : cache_data_798; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6957 = reset ? 185'h0 : cache_data_799; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6958 = reset ? 185'h0 : cache_data_800; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6959 = reset ? 185'h0 : cache_data_801; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6960 = reset ? 185'h0 : cache_data_802; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6961 = reset ? 185'h0 : cache_data_803; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6962 = reset ? 185'h0 : cache_data_804; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6963 = reset ? 185'h0 : cache_data_805; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6964 = reset ? 185'h0 : cache_data_806; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6965 = reset ? 185'h0 : cache_data_807; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6966 = reset ? 185'h0 : cache_data_808; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6967 = reset ? 185'h0 : cache_data_809; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6968 = reset ? 185'h0 : cache_data_810; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6969 = reset ? 185'h0 : cache_data_811; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6970 = reset ? 185'h0 : cache_data_812; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6971 = reset ? 185'h0 : cache_data_813; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6972 = reset ? 185'h0 : cache_data_814; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6973 = reset ? 185'h0 : cache_data_815; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6974 = reset ? 185'h0 : cache_data_816; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6975 = reset ? 185'h0 : cache_data_817; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6976 = reset ? 185'h0 : cache_data_818; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6977 = reset ? 185'h0 : cache_data_819; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6978 = reset ? 185'h0 : cache_data_820; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6979 = reset ? 185'h0 : cache_data_821; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6980 = reset ? 185'h0 : cache_data_822; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6981 = reset ? 185'h0 : cache_data_823; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6982 = reset ? 185'h0 : cache_data_824; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6983 = reset ? 185'h0 : cache_data_825; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6984 = reset ? 185'h0 : cache_data_826; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6985 = reset ? 185'h0 : cache_data_827; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6986 = reset ? 185'h0 : cache_data_828; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6987 = reset ? 185'h0 : cache_data_829; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6988 = reset ? 185'h0 : cache_data_830; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6989 = reset ? 185'h0 : cache_data_831; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6990 = reset ? 185'h0 : cache_data_832; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6991 = reset ? 185'h0 : cache_data_833; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6992 = reset ? 185'h0 : cache_data_834; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6993 = reset ? 185'h0 : cache_data_835; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6994 = reset ? 185'h0 : cache_data_836; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6995 = reset ? 185'h0 : cache_data_837; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6996 = reset ? 185'h0 : cache_data_838; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6997 = reset ? 185'h0 : cache_data_839; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6998 = reset ? 185'h0 : cache_data_840; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_6999 = reset ? 185'h0 : cache_data_841; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7000 = reset ? 185'h0 : cache_data_842; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7001 = reset ? 185'h0 : cache_data_843; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7002 = reset ? 185'h0 : cache_data_844; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7003 = reset ? 185'h0 : cache_data_845; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7004 = reset ? 185'h0 : cache_data_846; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7005 = reset ? 185'h0 : cache_data_847; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7006 = reset ? 185'h0 : cache_data_848; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7007 = reset ? 185'h0 : cache_data_849; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7008 = reset ? 185'h0 : cache_data_850; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7009 = reset ? 185'h0 : cache_data_851; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7010 = reset ? 185'h0 : cache_data_852; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7011 = reset ? 185'h0 : cache_data_853; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7012 = reset ? 185'h0 : cache_data_854; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7013 = reset ? 185'h0 : cache_data_855; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7014 = reset ? 185'h0 : cache_data_856; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7015 = reset ? 185'h0 : cache_data_857; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7016 = reset ? 185'h0 : cache_data_858; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7017 = reset ? 185'h0 : cache_data_859; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7018 = reset ? 185'h0 : cache_data_860; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7019 = reset ? 185'h0 : cache_data_861; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7020 = reset ? 185'h0 : cache_data_862; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7021 = reset ? 185'h0 : cache_data_863; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7022 = reset ? 185'h0 : cache_data_864; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7023 = reset ? 185'h0 : cache_data_865; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7024 = reset ? 185'h0 : cache_data_866; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7025 = reset ? 185'h0 : cache_data_867; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7026 = reset ? 185'h0 : cache_data_868; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7027 = reset ? 185'h0 : cache_data_869; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7028 = reset ? 185'h0 : cache_data_870; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7029 = reset ? 185'h0 : cache_data_871; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7030 = reset ? 185'h0 : cache_data_872; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7031 = reset ? 185'h0 : cache_data_873; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7032 = reset ? 185'h0 : cache_data_874; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7033 = reset ? 185'h0 : cache_data_875; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7034 = reset ? 185'h0 : cache_data_876; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7035 = reset ? 185'h0 : cache_data_877; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7036 = reset ? 185'h0 : cache_data_878; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7037 = reset ? 185'h0 : cache_data_879; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7038 = reset ? 185'h0 : cache_data_880; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7039 = reset ? 185'h0 : cache_data_881; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7040 = reset ? 185'h0 : cache_data_882; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7041 = reset ? 185'h0 : cache_data_883; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7042 = reset ? 185'h0 : cache_data_884; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7043 = reset ? 185'h0 : cache_data_885; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7044 = reset ? 185'h0 : cache_data_886; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7045 = reset ? 185'h0 : cache_data_887; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7046 = reset ? 185'h0 : cache_data_888; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7047 = reset ? 185'h0 : cache_data_889; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7048 = reset ? 185'h0 : cache_data_890; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7049 = reset ? 185'h0 : cache_data_891; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7050 = reset ? 185'h0 : cache_data_892; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7051 = reset ? 185'h0 : cache_data_893; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7052 = reset ? 185'h0 : cache_data_894; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7053 = reset ? 185'h0 : cache_data_895; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7054 = reset ? 185'h0 : cache_data_896; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7055 = reset ? 185'h0 : cache_data_897; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7056 = reset ? 185'h0 : cache_data_898; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7057 = reset ? 185'h0 : cache_data_899; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7058 = reset ? 185'h0 : cache_data_900; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7059 = reset ? 185'h0 : cache_data_901; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7060 = reset ? 185'h0 : cache_data_902; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7061 = reset ? 185'h0 : cache_data_903; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7062 = reset ? 185'h0 : cache_data_904; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7063 = reset ? 185'h0 : cache_data_905; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7064 = reset ? 185'h0 : cache_data_906; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7065 = reset ? 185'h0 : cache_data_907; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7066 = reset ? 185'h0 : cache_data_908; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7067 = reset ? 185'h0 : cache_data_909; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7068 = reset ? 185'h0 : cache_data_910; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7069 = reset ? 185'h0 : cache_data_911; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7070 = reset ? 185'h0 : cache_data_912; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7071 = reset ? 185'h0 : cache_data_913; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7072 = reset ? 185'h0 : cache_data_914; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7073 = reset ? 185'h0 : cache_data_915; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7074 = reset ? 185'h0 : cache_data_916; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7075 = reset ? 185'h0 : cache_data_917; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7076 = reset ? 185'h0 : cache_data_918; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7077 = reset ? 185'h0 : cache_data_919; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7078 = reset ? 185'h0 : cache_data_920; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7079 = reset ? 185'h0 : cache_data_921; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7080 = reset ? 185'h0 : cache_data_922; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7081 = reset ? 185'h0 : cache_data_923; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7082 = reset ? 185'h0 : cache_data_924; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7083 = reset ? 185'h0 : cache_data_925; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7084 = reset ? 185'h0 : cache_data_926; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7085 = reset ? 185'h0 : cache_data_927; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7086 = reset ? 185'h0 : cache_data_928; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7087 = reset ? 185'h0 : cache_data_929; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7088 = reset ? 185'h0 : cache_data_930; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7089 = reset ? 185'h0 : cache_data_931; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7090 = reset ? 185'h0 : cache_data_932; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7091 = reset ? 185'h0 : cache_data_933; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7092 = reset ? 185'h0 : cache_data_934; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7093 = reset ? 185'h0 : cache_data_935; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7094 = reset ? 185'h0 : cache_data_936; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7095 = reset ? 185'h0 : cache_data_937; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7096 = reset ? 185'h0 : cache_data_938; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7097 = reset ? 185'h0 : cache_data_939; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7098 = reset ? 185'h0 : cache_data_940; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7099 = reset ? 185'h0 : cache_data_941; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7100 = reset ? 185'h0 : cache_data_942; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7101 = reset ? 185'h0 : cache_data_943; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7102 = reset ? 185'h0 : cache_data_944; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7103 = reset ? 185'h0 : cache_data_945; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7104 = reset ? 185'h0 : cache_data_946; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7105 = reset ? 185'h0 : cache_data_947; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7106 = reset ? 185'h0 : cache_data_948; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7107 = reset ? 185'h0 : cache_data_949; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7108 = reset ? 185'h0 : cache_data_950; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7109 = reset ? 185'h0 : cache_data_951; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7110 = reset ? 185'h0 : cache_data_952; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7111 = reset ? 185'h0 : cache_data_953; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7112 = reset ? 185'h0 : cache_data_954; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7113 = reset ? 185'h0 : cache_data_955; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7114 = reset ? 185'h0 : cache_data_956; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7115 = reset ? 185'h0 : cache_data_957; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7116 = reset ? 185'h0 : cache_data_958; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7117 = reset ? 185'h0 : cache_data_959; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7118 = reset ? 185'h0 : cache_data_960; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7119 = reset ? 185'h0 : cache_data_961; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7120 = reset ? 185'h0 : cache_data_962; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7121 = reset ? 185'h0 : cache_data_963; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7122 = reset ? 185'h0 : cache_data_964; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7123 = reset ? 185'h0 : cache_data_965; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7124 = reset ? 185'h0 : cache_data_966; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7125 = reset ? 185'h0 : cache_data_967; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7126 = reset ? 185'h0 : cache_data_968; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7127 = reset ? 185'h0 : cache_data_969; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7128 = reset ? 185'h0 : cache_data_970; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7129 = reset ? 185'h0 : cache_data_971; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7130 = reset ? 185'h0 : cache_data_972; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7131 = reset ? 185'h0 : cache_data_973; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7132 = reset ? 185'h0 : cache_data_974; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7133 = reset ? 185'h0 : cache_data_975; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7134 = reset ? 185'h0 : cache_data_976; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7135 = reset ? 185'h0 : cache_data_977; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7136 = reset ? 185'h0 : cache_data_978; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7137 = reset ? 185'h0 : cache_data_979; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7138 = reset ? 185'h0 : cache_data_980; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7139 = reset ? 185'h0 : cache_data_981; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7140 = reset ? 185'h0 : cache_data_982; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7141 = reset ? 185'h0 : cache_data_983; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7142 = reset ? 185'h0 : cache_data_984; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7143 = reset ? 185'h0 : cache_data_985; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7144 = reset ? 185'h0 : cache_data_986; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7145 = reset ? 185'h0 : cache_data_987; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7146 = reset ? 185'h0 : cache_data_988; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7147 = reset ? 185'h0 : cache_data_989; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7148 = reset ? 185'h0 : cache_data_990; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7149 = reset ? 185'h0 : cache_data_991; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7150 = reset ? 185'h0 : cache_data_992; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7151 = reset ? 185'h0 : cache_data_993; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7152 = reset ? 185'h0 : cache_data_994; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7153 = reset ? 185'h0 : cache_data_995; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7154 = reset ? 185'h0 : cache_data_996; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7155 = reset ? 185'h0 : cache_data_997; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7156 = reset ? 185'h0 : cache_data_998; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7157 = reset ? 185'h0 : cache_data_999; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7158 = reset ? 185'h0 : cache_data_1000; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7159 = reset ? 185'h0 : cache_data_1001; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7160 = reset ? 185'h0 : cache_data_1002; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7161 = reset ? 185'h0 : cache_data_1003; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7162 = reset ? 185'h0 : cache_data_1004; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7163 = reset ? 185'h0 : cache_data_1005; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7164 = reset ? 185'h0 : cache_data_1006; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7165 = reset ? 185'h0 : cache_data_1007; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7166 = reset ? 185'h0 : cache_data_1008; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7167 = reset ? 185'h0 : cache_data_1009; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7168 = reset ? 185'h0 : cache_data_1010; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7169 = reset ? 185'h0 : cache_data_1011; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7170 = reset ? 185'h0 : cache_data_1012; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7171 = reset ? 185'h0 : cache_data_1013; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7172 = reset ? 185'h0 : cache_data_1014; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7173 = reset ? 185'h0 : cache_data_1015; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7174 = reset ? 185'h0 : cache_data_1016; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7175 = reset ? 185'h0 : cache_data_1017; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7176 = reset ? 185'h0 : cache_data_1018; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7177 = reset ? 185'h0 : cache_data_1019; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7178 = reset ? 185'h0 : cache_data_1020; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7179 = reset ? 185'h0 : cache_data_1021; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7180 = reset ? 185'h0 : cache_data_1022; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _GEN_7181 = reset ? 185'h0 : cache_data_1023; // @[icache.scala 128:24 131:21 47:23]
  wire [184:0] _cache_data_T_6 = {_GEN_4095[184],1'h0,_GEN_4095[182:0]}; // @[Cat.scala 31:58]
  wire [184:0] _GEN_9230 = 10'h0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6158; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9231 = 10'h1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6159; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9232 = 10'h2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6160; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9233 = 10'h3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6161; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9234 = 10'h4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6162; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9235 = 10'h5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6163; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9236 = 10'h6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6164; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9237 = 10'h7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6165; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9238 = 10'h8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6166; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9239 = 10'h9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6167; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9240 = 10'ha == _dirty_T_1 ? _cache_data_T_6 : _GEN_6168; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9241 = 10'hb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6169; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9242 = 10'hc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6170; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9243 = 10'hd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6171; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9244 = 10'he == _dirty_T_1 ? _cache_data_T_6 : _GEN_6172; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9245 = 10'hf == _dirty_T_1 ? _cache_data_T_6 : _GEN_6173; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9246 = 10'h10 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6174; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9247 = 10'h11 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6175; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9248 = 10'h12 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6176; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9249 = 10'h13 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6177; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9250 = 10'h14 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6178; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9251 = 10'h15 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6179; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9252 = 10'h16 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6180; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9253 = 10'h17 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6181; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9254 = 10'h18 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6182; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9255 = 10'h19 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6183; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9256 = 10'h1a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6184; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9257 = 10'h1b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6185; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9258 = 10'h1c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6186; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9259 = 10'h1d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6187; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9260 = 10'h1e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6188; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9261 = 10'h1f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6189; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9262 = 10'h20 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6190; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9263 = 10'h21 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6191; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9264 = 10'h22 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6192; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9265 = 10'h23 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6193; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9266 = 10'h24 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6194; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9267 = 10'h25 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6195; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9268 = 10'h26 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6196; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9269 = 10'h27 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6197; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9270 = 10'h28 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6198; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9271 = 10'h29 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6199; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9272 = 10'h2a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6200; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9273 = 10'h2b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6201; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9274 = 10'h2c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6202; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9275 = 10'h2d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6203; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9276 = 10'h2e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6204; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9277 = 10'h2f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6205; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9278 = 10'h30 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6206; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9279 = 10'h31 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6207; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9280 = 10'h32 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6208; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9281 = 10'h33 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6209; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9282 = 10'h34 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6210; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9283 = 10'h35 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6211; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9284 = 10'h36 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6212; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9285 = 10'h37 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6213; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9286 = 10'h38 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6214; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9287 = 10'h39 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6215; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9288 = 10'h3a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6216; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9289 = 10'h3b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6217; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9290 = 10'h3c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6218; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9291 = 10'h3d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6219; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9292 = 10'h3e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6220; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9293 = 10'h3f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6221; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9294 = 10'h40 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6222; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9295 = 10'h41 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6223; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9296 = 10'h42 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6224; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9297 = 10'h43 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6225; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9298 = 10'h44 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6226; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9299 = 10'h45 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6227; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9300 = 10'h46 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6228; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9301 = 10'h47 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6229; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9302 = 10'h48 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6230; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9303 = 10'h49 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6231; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9304 = 10'h4a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6232; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9305 = 10'h4b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6233; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9306 = 10'h4c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6234; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9307 = 10'h4d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6235; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9308 = 10'h4e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6236; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9309 = 10'h4f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6237; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9310 = 10'h50 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6238; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9311 = 10'h51 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6239; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9312 = 10'h52 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6240; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9313 = 10'h53 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6241; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9314 = 10'h54 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6242; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9315 = 10'h55 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6243; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9316 = 10'h56 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6244; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9317 = 10'h57 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6245; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9318 = 10'h58 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6246; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9319 = 10'h59 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6247; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9320 = 10'h5a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6248; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9321 = 10'h5b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6249; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9322 = 10'h5c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6250; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9323 = 10'h5d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6251; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9324 = 10'h5e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6252; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9325 = 10'h5f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6253; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9326 = 10'h60 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6254; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9327 = 10'h61 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6255; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9328 = 10'h62 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6256; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9329 = 10'h63 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6257; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9330 = 10'h64 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6258; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9331 = 10'h65 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6259; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9332 = 10'h66 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6260; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9333 = 10'h67 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6261; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9334 = 10'h68 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6262; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9335 = 10'h69 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6263; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9336 = 10'h6a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6264; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9337 = 10'h6b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6265; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9338 = 10'h6c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6266; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9339 = 10'h6d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6267; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9340 = 10'h6e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6268; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9341 = 10'h6f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6269; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9342 = 10'h70 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6270; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9343 = 10'h71 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6271; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9344 = 10'h72 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6272; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9345 = 10'h73 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6273; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9346 = 10'h74 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6274; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9347 = 10'h75 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6275; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9348 = 10'h76 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6276; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9349 = 10'h77 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6277; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9350 = 10'h78 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6278; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9351 = 10'h79 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6279; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9352 = 10'h7a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6280; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9353 = 10'h7b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6281; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9354 = 10'h7c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6282; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9355 = 10'h7d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6283; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9356 = 10'h7e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6284; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9357 = 10'h7f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6285; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9358 = 10'h80 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6286; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9359 = 10'h81 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6287; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9360 = 10'h82 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6288; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9361 = 10'h83 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6289; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9362 = 10'h84 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6290; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9363 = 10'h85 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6291; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9364 = 10'h86 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6292; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9365 = 10'h87 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6293; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9366 = 10'h88 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6294; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9367 = 10'h89 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6295; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9368 = 10'h8a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6296; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9369 = 10'h8b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6297; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9370 = 10'h8c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6298; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9371 = 10'h8d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6299; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9372 = 10'h8e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6300; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9373 = 10'h8f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6301; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9374 = 10'h90 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6302; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9375 = 10'h91 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6303; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9376 = 10'h92 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6304; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9377 = 10'h93 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6305; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9378 = 10'h94 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6306; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9379 = 10'h95 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6307; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9380 = 10'h96 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6308; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9381 = 10'h97 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6309; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9382 = 10'h98 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6310; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9383 = 10'h99 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6311; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9384 = 10'h9a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6312; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9385 = 10'h9b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6313; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9386 = 10'h9c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6314; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9387 = 10'h9d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6315; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9388 = 10'h9e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6316; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9389 = 10'h9f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6317; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9390 = 10'ha0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6318; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9391 = 10'ha1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6319; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9392 = 10'ha2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6320; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9393 = 10'ha3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6321; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9394 = 10'ha4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6322; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9395 = 10'ha5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6323; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9396 = 10'ha6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6324; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9397 = 10'ha7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6325; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9398 = 10'ha8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6326; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9399 = 10'ha9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6327; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9400 = 10'haa == _dirty_T_1 ? _cache_data_T_6 : _GEN_6328; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9401 = 10'hab == _dirty_T_1 ? _cache_data_T_6 : _GEN_6329; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9402 = 10'hac == _dirty_T_1 ? _cache_data_T_6 : _GEN_6330; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9403 = 10'had == _dirty_T_1 ? _cache_data_T_6 : _GEN_6331; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9404 = 10'hae == _dirty_T_1 ? _cache_data_T_6 : _GEN_6332; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9405 = 10'haf == _dirty_T_1 ? _cache_data_T_6 : _GEN_6333; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9406 = 10'hb0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6334; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9407 = 10'hb1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6335; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9408 = 10'hb2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6336; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9409 = 10'hb3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6337; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9410 = 10'hb4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6338; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9411 = 10'hb5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6339; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9412 = 10'hb6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6340; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9413 = 10'hb7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6341; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9414 = 10'hb8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6342; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9415 = 10'hb9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6343; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9416 = 10'hba == _dirty_T_1 ? _cache_data_T_6 : _GEN_6344; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9417 = 10'hbb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6345; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9418 = 10'hbc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6346; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9419 = 10'hbd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6347; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9420 = 10'hbe == _dirty_T_1 ? _cache_data_T_6 : _GEN_6348; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9421 = 10'hbf == _dirty_T_1 ? _cache_data_T_6 : _GEN_6349; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9422 = 10'hc0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6350; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9423 = 10'hc1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6351; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9424 = 10'hc2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6352; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9425 = 10'hc3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6353; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9426 = 10'hc4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6354; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9427 = 10'hc5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6355; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9428 = 10'hc6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6356; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9429 = 10'hc7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6357; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9430 = 10'hc8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6358; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9431 = 10'hc9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6359; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9432 = 10'hca == _dirty_T_1 ? _cache_data_T_6 : _GEN_6360; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9433 = 10'hcb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6361; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9434 = 10'hcc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6362; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9435 = 10'hcd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6363; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9436 = 10'hce == _dirty_T_1 ? _cache_data_T_6 : _GEN_6364; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9437 = 10'hcf == _dirty_T_1 ? _cache_data_T_6 : _GEN_6365; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9438 = 10'hd0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6366; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9439 = 10'hd1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6367; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9440 = 10'hd2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6368; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9441 = 10'hd3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6369; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9442 = 10'hd4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6370; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9443 = 10'hd5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6371; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9444 = 10'hd6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6372; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9445 = 10'hd7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6373; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9446 = 10'hd8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6374; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9447 = 10'hd9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6375; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9448 = 10'hda == _dirty_T_1 ? _cache_data_T_6 : _GEN_6376; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9449 = 10'hdb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6377; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9450 = 10'hdc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6378; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9451 = 10'hdd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6379; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9452 = 10'hde == _dirty_T_1 ? _cache_data_T_6 : _GEN_6380; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9453 = 10'hdf == _dirty_T_1 ? _cache_data_T_6 : _GEN_6381; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9454 = 10'he0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6382; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9455 = 10'he1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6383; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9456 = 10'he2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6384; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9457 = 10'he3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6385; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9458 = 10'he4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6386; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9459 = 10'he5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6387; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9460 = 10'he6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6388; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9461 = 10'he7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6389; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9462 = 10'he8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6390; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9463 = 10'he9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6391; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9464 = 10'hea == _dirty_T_1 ? _cache_data_T_6 : _GEN_6392; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9465 = 10'heb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6393; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9466 = 10'hec == _dirty_T_1 ? _cache_data_T_6 : _GEN_6394; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9467 = 10'hed == _dirty_T_1 ? _cache_data_T_6 : _GEN_6395; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9468 = 10'hee == _dirty_T_1 ? _cache_data_T_6 : _GEN_6396; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9469 = 10'hef == _dirty_T_1 ? _cache_data_T_6 : _GEN_6397; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9470 = 10'hf0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6398; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9471 = 10'hf1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6399; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9472 = 10'hf2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6400; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9473 = 10'hf3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6401; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9474 = 10'hf4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6402; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9475 = 10'hf5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6403; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9476 = 10'hf6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6404; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9477 = 10'hf7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6405; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9478 = 10'hf8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6406; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9479 = 10'hf9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6407; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9480 = 10'hfa == _dirty_T_1 ? _cache_data_T_6 : _GEN_6408; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9481 = 10'hfb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6409; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9482 = 10'hfc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6410; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9483 = 10'hfd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6411; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9484 = 10'hfe == _dirty_T_1 ? _cache_data_T_6 : _GEN_6412; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9485 = 10'hff == _dirty_T_1 ? _cache_data_T_6 : _GEN_6413; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9486 = 10'h100 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6414; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9487 = 10'h101 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6415; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9488 = 10'h102 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6416; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9489 = 10'h103 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6417; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9490 = 10'h104 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6418; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9491 = 10'h105 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6419; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9492 = 10'h106 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6420; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9493 = 10'h107 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6421; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9494 = 10'h108 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6422; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9495 = 10'h109 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6423; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9496 = 10'h10a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6424; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9497 = 10'h10b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6425; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9498 = 10'h10c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6426; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9499 = 10'h10d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6427; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9500 = 10'h10e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6428; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9501 = 10'h10f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6429; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9502 = 10'h110 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6430; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9503 = 10'h111 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6431; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9504 = 10'h112 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6432; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9505 = 10'h113 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6433; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9506 = 10'h114 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6434; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9507 = 10'h115 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6435; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9508 = 10'h116 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6436; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9509 = 10'h117 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6437; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9510 = 10'h118 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6438; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9511 = 10'h119 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6439; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9512 = 10'h11a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6440; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9513 = 10'h11b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6441; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9514 = 10'h11c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6442; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9515 = 10'h11d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6443; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9516 = 10'h11e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6444; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9517 = 10'h11f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6445; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9518 = 10'h120 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6446; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9519 = 10'h121 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6447; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9520 = 10'h122 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6448; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9521 = 10'h123 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6449; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9522 = 10'h124 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6450; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9523 = 10'h125 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6451; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9524 = 10'h126 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6452; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9525 = 10'h127 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6453; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9526 = 10'h128 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6454; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9527 = 10'h129 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6455; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9528 = 10'h12a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6456; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9529 = 10'h12b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6457; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9530 = 10'h12c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6458; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9531 = 10'h12d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6459; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9532 = 10'h12e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6460; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9533 = 10'h12f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6461; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9534 = 10'h130 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6462; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9535 = 10'h131 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6463; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9536 = 10'h132 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6464; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9537 = 10'h133 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6465; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9538 = 10'h134 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6466; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9539 = 10'h135 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6467; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9540 = 10'h136 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6468; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9541 = 10'h137 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6469; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9542 = 10'h138 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6470; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9543 = 10'h139 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6471; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9544 = 10'h13a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6472; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9545 = 10'h13b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6473; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9546 = 10'h13c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6474; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9547 = 10'h13d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6475; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9548 = 10'h13e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6476; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9549 = 10'h13f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6477; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9550 = 10'h140 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6478; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9551 = 10'h141 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6479; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9552 = 10'h142 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6480; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9553 = 10'h143 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6481; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9554 = 10'h144 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6482; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9555 = 10'h145 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6483; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9556 = 10'h146 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6484; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9557 = 10'h147 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6485; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9558 = 10'h148 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6486; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9559 = 10'h149 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6487; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9560 = 10'h14a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6488; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9561 = 10'h14b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6489; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9562 = 10'h14c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6490; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9563 = 10'h14d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6491; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9564 = 10'h14e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6492; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9565 = 10'h14f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6493; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9566 = 10'h150 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6494; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9567 = 10'h151 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6495; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9568 = 10'h152 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6496; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9569 = 10'h153 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6497; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9570 = 10'h154 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6498; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9571 = 10'h155 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6499; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9572 = 10'h156 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6500; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9573 = 10'h157 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6501; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9574 = 10'h158 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6502; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9575 = 10'h159 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6503; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9576 = 10'h15a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6504; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9577 = 10'h15b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6505; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9578 = 10'h15c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6506; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9579 = 10'h15d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6507; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9580 = 10'h15e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6508; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9581 = 10'h15f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6509; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9582 = 10'h160 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6510; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9583 = 10'h161 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6511; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9584 = 10'h162 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6512; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9585 = 10'h163 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6513; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9586 = 10'h164 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6514; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9587 = 10'h165 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6515; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9588 = 10'h166 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6516; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9589 = 10'h167 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6517; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9590 = 10'h168 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6518; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9591 = 10'h169 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6519; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9592 = 10'h16a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6520; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9593 = 10'h16b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6521; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9594 = 10'h16c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6522; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9595 = 10'h16d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6523; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9596 = 10'h16e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6524; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9597 = 10'h16f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6525; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9598 = 10'h170 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6526; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9599 = 10'h171 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6527; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9600 = 10'h172 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6528; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9601 = 10'h173 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6529; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9602 = 10'h174 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6530; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9603 = 10'h175 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6531; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9604 = 10'h176 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6532; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9605 = 10'h177 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6533; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9606 = 10'h178 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6534; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9607 = 10'h179 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6535; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9608 = 10'h17a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6536; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9609 = 10'h17b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6537; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9610 = 10'h17c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6538; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9611 = 10'h17d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6539; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9612 = 10'h17e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6540; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9613 = 10'h17f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6541; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9614 = 10'h180 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6542; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9615 = 10'h181 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6543; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9616 = 10'h182 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6544; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9617 = 10'h183 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6545; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9618 = 10'h184 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6546; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9619 = 10'h185 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6547; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9620 = 10'h186 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6548; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9621 = 10'h187 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6549; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9622 = 10'h188 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6550; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9623 = 10'h189 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6551; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9624 = 10'h18a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6552; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9625 = 10'h18b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6553; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9626 = 10'h18c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6554; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9627 = 10'h18d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6555; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9628 = 10'h18e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6556; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9629 = 10'h18f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6557; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9630 = 10'h190 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6558; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9631 = 10'h191 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6559; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9632 = 10'h192 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6560; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9633 = 10'h193 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6561; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9634 = 10'h194 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6562; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9635 = 10'h195 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6563; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9636 = 10'h196 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6564; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9637 = 10'h197 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6565; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9638 = 10'h198 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6566; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9639 = 10'h199 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6567; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9640 = 10'h19a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6568; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9641 = 10'h19b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6569; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9642 = 10'h19c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6570; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9643 = 10'h19d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6571; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9644 = 10'h19e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6572; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9645 = 10'h19f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6573; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9646 = 10'h1a0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6574; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9647 = 10'h1a1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6575; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9648 = 10'h1a2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6576; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9649 = 10'h1a3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6577; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9650 = 10'h1a4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6578; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9651 = 10'h1a5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6579; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9652 = 10'h1a6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6580; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9653 = 10'h1a7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6581; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9654 = 10'h1a8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6582; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9655 = 10'h1a9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6583; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9656 = 10'h1aa == _dirty_T_1 ? _cache_data_T_6 : _GEN_6584; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9657 = 10'h1ab == _dirty_T_1 ? _cache_data_T_6 : _GEN_6585; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9658 = 10'h1ac == _dirty_T_1 ? _cache_data_T_6 : _GEN_6586; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9659 = 10'h1ad == _dirty_T_1 ? _cache_data_T_6 : _GEN_6587; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9660 = 10'h1ae == _dirty_T_1 ? _cache_data_T_6 : _GEN_6588; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9661 = 10'h1af == _dirty_T_1 ? _cache_data_T_6 : _GEN_6589; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9662 = 10'h1b0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6590; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9663 = 10'h1b1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6591; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9664 = 10'h1b2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6592; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9665 = 10'h1b3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6593; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9666 = 10'h1b4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6594; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9667 = 10'h1b5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6595; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9668 = 10'h1b6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6596; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9669 = 10'h1b7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6597; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9670 = 10'h1b8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6598; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9671 = 10'h1b9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6599; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9672 = 10'h1ba == _dirty_T_1 ? _cache_data_T_6 : _GEN_6600; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9673 = 10'h1bb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6601; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9674 = 10'h1bc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6602; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9675 = 10'h1bd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6603; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9676 = 10'h1be == _dirty_T_1 ? _cache_data_T_6 : _GEN_6604; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9677 = 10'h1bf == _dirty_T_1 ? _cache_data_T_6 : _GEN_6605; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9678 = 10'h1c0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6606; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9679 = 10'h1c1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6607; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9680 = 10'h1c2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6608; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9681 = 10'h1c3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6609; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9682 = 10'h1c4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6610; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9683 = 10'h1c5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6611; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9684 = 10'h1c6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6612; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9685 = 10'h1c7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6613; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9686 = 10'h1c8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6614; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9687 = 10'h1c9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6615; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9688 = 10'h1ca == _dirty_T_1 ? _cache_data_T_6 : _GEN_6616; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9689 = 10'h1cb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6617; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9690 = 10'h1cc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6618; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9691 = 10'h1cd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6619; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9692 = 10'h1ce == _dirty_T_1 ? _cache_data_T_6 : _GEN_6620; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9693 = 10'h1cf == _dirty_T_1 ? _cache_data_T_6 : _GEN_6621; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9694 = 10'h1d0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6622; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9695 = 10'h1d1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6623; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9696 = 10'h1d2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6624; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9697 = 10'h1d3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6625; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9698 = 10'h1d4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6626; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9699 = 10'h1d5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6627; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9700 = 10'h1d6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6628; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9701 = 10'h1d7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6629; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9702 = 10'h1d8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6630; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9703 = 10'h1d9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6631; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9704 = 10'h1da == _dirty_T_1 ? _cache_data_T_6 : _GEN_6632; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9705 = 10'h1db == _dirty_T_1 ? _cache_data_T_6 : _GEN_6633; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9706 = 10'h1dc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6634; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9707 = 10'h1dd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6635; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9708 = 10'h1de == _dirty_T_1 ? _cache_data_T_6 : _GEN_6636; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9709 = 10'h1df == _dirty_T_1 ? _cache_data_T_6 : _GEN_6637; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9710 = 10'h1e0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6638; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9711 = 10'h1e1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6639; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9712 = 10'h1e2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6640; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9713 = 10'h1e3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6641; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9714 = 10'h1e4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6642; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9715 = 10'h1e5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6643; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9716 = 10'h1e6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6644; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9717 = 10'h1e7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6645; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9718 = 10'h1e8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6646; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9719 = 10'h1e9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6647; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9720 = 10'h1ea == _dirty_T_1 ? _cache_data_T_6 : _GEN_6648; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9721 = 10'h1eb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6649; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9722 = 10'h1ec == _dirty_T_1 ? _cache_data_T_6 : _GEN_6650; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9723 = 10'h1ed == _dirty_T_1 ? _cache_data_T_6 : _GEN_6651; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9724 = 10'h1ee == _dirty_T_1 ? _cache_data_T_6 : _GEN_6652; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9725 = 10'h1ef == _dirty_T_1 ? _cache_data_T_6 : _GEN_6653; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9726 = 10'h1f0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6654; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9727 = 10'h1f1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6655; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9728 = 10'h1f2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6656; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9729 = 10'h1f3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6657; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9730 = 10'h1f4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6658; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9731 = 10'h1f5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6659; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9732 = 10'h1f6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6660; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9733 = 10'h1f7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6661; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9734 = 10'h1f8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6662; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9735 = 10'h1f9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6663; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9736 = 10'h1fa == _dirty_T_1 ? _cache_data_T_6 : _GEN_6664; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9737 = 10'h1fb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6665; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9738 = 10'h1fc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6666; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9739 = 10'h1fd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6667; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9740 = 10'h1fe == _dirty_T_1 ? _cache_data_T_6 : _GEN_6668; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9741 = 10'h1ff == _dirty_T_1 ? _cache_data_T_6 : _GEN_6669; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9742 = 10'h200 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6670; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9743 = 10'h201 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6671; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9744 = 10'h202 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6672; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9745 = 10'h203 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6673; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9746 = 10'h204 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6674; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9747 = 10'h205 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6675; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9748 = 10'h206 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6676; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9749 = 10'h207 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6677; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9750 = 10'h208 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6678; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9751 = 10'h209 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6679; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9752 = 10'h20a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6680; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9753 = 10'h20b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6681; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9754 = 10'h20c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6682; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9755 = 10'h20d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6683; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9756 = 10'h20e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6684; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9757 = 10'h20f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6685; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9758 = 10'h210 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6686; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9759 = 10'h211 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6687; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9760 = 10'h212 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6688; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9761 = 10'h213 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6689; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9762 = 10'h214 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6690; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9763 = 10'h215 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6691; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9764 = 10'h216 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6692; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9765 = 10'h217 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6693; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9766 = 10'h218 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6694; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9767 = 10'h219 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6695; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9768 = 10'h21a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6696; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9769 = 10'h21b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6697; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9770 = 10'h21c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6698; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9771 = 10'h21d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6699; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9772 = 10'h21e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6700; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9773 = 10'h21f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6701; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9774 = 10'h220 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6702; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9775 = 10'h221 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6703; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9776 = 10'h222 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6704; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9777 = 10'h223 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6705; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9778 = 10'h224 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6706; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9779 = 10'h225 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6707; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9780 = 10'h226 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6708; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9781 = 10'h227 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6709; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9782 = 10'h228 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6710; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9783 = 10'h229 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6711; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9784 = 10'h22a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6712; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9785 = 10'h22b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6713; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9786 = 10'h22c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6714; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9787 = 10'h22d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6715; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9788 = 10'h22e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6716; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9789 = 10'h22f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6717; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9790 = 10'h230 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6718; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9791 = 10'h231 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6719; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9792 = 10'h232 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6720; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9793 = 10'h233 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6721; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9794 = 10'h234 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6722; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9795 = 10'h235 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6723; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9796 = 10'h236 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6724; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9797 = 10'h237 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6725; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9798 = 10'h238 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6726; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9799 = 10'h239 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6727; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9800 = 10'h23a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6728; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9801 = 10'h23b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6729; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9802 = 10'h23c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6730; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9803 = 10'h23d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6731; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9804 = 10'h23e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6732; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9805 = 10'h23f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6733; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9806 = 10'h240 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6734; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9807 = 10'h241 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6735; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9808 = 10'h242 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6736; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9809 = 10'h243 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6737; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9810 = 10'h244 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6738; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9811 = 10'h245 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6739; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9812 = 10'h246 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6740; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9813 = 10'h247 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6741; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9814 = 10'h248 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6742; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9815 = 10'h249 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6743; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9816 = 10'h24a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6744; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9817 = 10'h24b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6745; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9818 = 10'h24c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6746; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9819 = 10'h24d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6747; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9820 = 10'h24e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6748; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9821 = 10'h24f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6749; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9822 = 10'h250 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6750; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9823 = 10'h251 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6751; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9824 = 10'h252 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6752; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9825 = 10'h253 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6753; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9826 = 10'h254 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6754; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9827 = 10'h255 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6755; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9828 = 10'h256 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6756; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9829 = 10'h257 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6757; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9830 = 10'h258 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6758; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9831 = 10'h259 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6759; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9832 = 10'h25a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6760; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9833 = 10'h25b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6761; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9834 = 10'h25c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6762; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9835 = 10'h25d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6763; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9836 = 10'h25e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6764; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9837 = 10'h25f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6765; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9838 = 10'h260 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6766; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9839 = 10'h261 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6767; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9840 = 10'h262 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6768; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9841 = 10'h263 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6769; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9842 = 10'h264 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6770; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9843 = 10'h265 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6771; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9844 = 10'h266 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6772; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9845 = 10'h267 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6773; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9846 = 10'h268 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6774; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9847 = 10'h269 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6775; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9848 = 10'h26a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6776; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9849 = 10'h26b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6777; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9850 = 10'h26c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6778; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9851 = 10'h26d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6779; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9852 = 10'h26e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6780; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9853 = 10'h26f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6781; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9854 = 10'h270 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6782; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9855 = 10'h271 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6783; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9856 = 10'h272 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6784; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9857 = 10'h273 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6785; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9858 = 10'h274 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6786; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9859 = 10'h275 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6787; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9860 = 10'h276 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6788; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9861 = 10'h277 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6789; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9862 = 10'h278 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6790; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9863 = 10'h279 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6791; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9864 = 10'h27a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6792; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9865 = 10'h27b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6793; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9866 = 10'h27c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6794; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9867 = 10'h27d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6795; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9868 = 10'h27e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6796; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9869 = 10'h27f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6797; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9870 = 10'h280 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6798; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9871 = 10'h281 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6799; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9872 = 10'h282 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6800; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9873 = 10'h283 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6801; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9874 = 10'h284 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6802; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9875 = 10'h285 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6803; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9876 = 10'h286 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6804; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9877 = 10'h287 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6805; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9878 = 10'h288 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6806; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9879 = 10'h289 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6807; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9880 = 10'h28a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6808; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9881 = 10'h28b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6809; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9882 = 10'h28c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6810; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9883 = 10'h28d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6811; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9884 = 10'h28e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6812; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9885 = 10'h28f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6813; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9886 = 10'h290 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6814; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9887 = 10'h291 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6815; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9888 = 10'h292 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6816; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9889 = 10'h293 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6817; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9890 = 10'h294 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6818; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9891 = 10'h295 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6819; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9892 = 10'h296 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6820; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9893 = 10'h297 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6821; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9894 = 10'h298 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6822; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9895 = 10'h299 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6823; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9896 = 10'h29a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6824; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9897 = 10'h29b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6825; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9898 = 10'h29c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6826; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9899 = 10'h29d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6827; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9900 = 10'h29e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6828; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9901 = 10'h29f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6829; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9902 = 10'h2a0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6830; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9903 = 10'h2a1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6831; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9904 = 10'h2a2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6832; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9905 = 10'h2a3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6833; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9906 = 10'h2a4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6834; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9907 = 10'h2a5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6835; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9908 = 10'h2a6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6836; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9909 = 10'h2a7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6837; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9910 = 10'h2a8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6838; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9911 = 10'h2a9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6839; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9912 = 10'h2aa == _dirty_T_1 ? _cache_data_T_6 : _GEN_6840; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9913 = 10'h2ab == _dirty_T_1 ? _cache_data_T_6 : _GEN_6841; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9914 = 10'h2ac == _dirty_T_1 ? _cache_data_T_6 : _GEN_6842; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9915 = 10'h2ad == _dirty_T_1 ? _cache_data_T_6 : _GEN_6843; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9916 = 10'h2ae == _dirty_T_1 ? _cache_data_T_6 : _GEN_6844; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9917 = 10'h2af == _dirty_T_1 ? _cache_data_T_6 : _GEN_6845; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9918 = 10'h2b0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6846; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9919 = 10'h2b1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6847; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9920 = 10'h2b2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6848; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9921 = 10'h2b3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6849; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9922 = 10'h2b4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6850; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9923 = 10'h2b5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6851; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9924 = 10'h2b6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6852; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9925 = 10'h2b7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6853; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9926 = 10'h2b8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6854; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9927 = 10'h2b9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6855; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9928 = 10'h2ba == _dirty_T_1 ? _cache_data_T_6 : _GEN_6856; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9929 = 10'h2bb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6857; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9930 = 10'h2bc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6858; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9931 = 10'h2bd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6859; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9932 = 10'h2be == _dirty_T_1 ? _cache_data_T_6 : _GEN_6860; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9933 = 10'h2bf == _dirty_T_1 ? _cache_data_T_6 : _GEN_6861; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9934 = 10'h2c0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6862; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9935 = 10'h2c1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6863; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9936 = 10'h2c2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6864; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9937 = 10'h2c3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6865; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9938 = 10'h2c4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6866; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9939 = 10'h2c5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6867; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9940 = 10'h2c6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6868; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9941 = 10'h2c7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6869; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9942 = 10'h2c8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6870; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9943 = 10'h2c9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6871; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9944 = 10'h2ca == _dirty_T_1 ? _cache_data_T_6 : _GEN_6872; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9945 = 10'h2cb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6873; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9946 = 10'h2cc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6874; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9947 = 10'h2cd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6875; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9948 = 10'h2ce == _dirty_T_1 ? _cache_data_T_6 : _GEN_6876; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9949 = 10'h2cf == _dirty_T_1 ? _cache_data_T_6 : _GEN_6877; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9950 = 10'h2d0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6878; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9951 = 10'h2d1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6879; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9952 = 10'h2d2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6880; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9953 = 10'h2d3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6881; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9954 = 10'h2d4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6882; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9955 = 10'h2d5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6883; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9956 = 10'h2d6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6884; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9957 = 10'h2d7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6885; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9958 = 10'h2d8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6886; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9959 = 10'h2d9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6887; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9960 = 10'h2da == _dirty_T_1 ? _cache_data_T_6 : _GEN_6888; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9961 = 10'h2db == _dirty_T_1 ? _cache_data_T_6 : _GEN_6889; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9962 = 10'h2dc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6890; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9963 = 10'h2dd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6891; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9964 = 10'h2de == _dirty_T_1 ? _cache_data_T_6 : _GEN_6892; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9965 = 10'h2df == _dirty_T_1 ? _cache_data_T_6 : _GEN_6893; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9966 = 10'h2e0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6894; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9967 = 10'h2e1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6895; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9968 = 10'h2e2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6896; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9969 = 10'h2e3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6897; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9970 = 10'h2e4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6898; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9971 = 10'h2e5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6899; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9972 = 10'h2e6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6900; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9973 = 10'h2e7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6901; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9974 = 10'h2e8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6902; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9975 = 10'h2e9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6903; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9976 = 10'h2ea == _dirty_T_1 ? _cache_data_T_6 : _GEN_6904; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9977 = 10'h2eb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6905; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9978 = 10'h2ec == _dirty_T_1 ? _cache_data_T_6 : _GEN_6906; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9979 = 10'h2ed == _dirty_T_1 ? _cache_data_T_6 : _GEN_6907; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9980 = 10'h2ee == _dirty_T_1 ? _cache_data_T_6 : _GEN_6908; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9981 = 10'h2ef == _dirty_T_1 ? _cache_data_T_6 : _GEN_6909; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9982 = 10'h2f0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6910; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9983 = 10'h2f1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6911; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9984 = 10'h2f2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6912; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9985 = 10'h2f3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6913; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9986 = 10'h2f4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6914; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9987 = 10'h2f5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6915; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9988 = 10'h2f6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6916; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9989 = 10'h2f7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6917; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9990 = 10'h2f8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6918; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9991 = 10'h2f9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6919; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9992 = 10'h2fa == _dirty_T_1 ? _cache_data_T_6 : _GEN_6920; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9993 = 10'h2fb == _dirty_T_1 ? _cache_data_T_6 : _GEN_6921; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9994 = 10'h2fc == _dirty_T_1 ? _cache_data_T_6 : _GEN_6922; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9995 = 10'h2fd == _dirty_T_1 ? _cache_data_T_6 : _GEN_6923; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9996 = 10'h2fe == _dirty_T_1 ? _cache_data_T_6 : _GEN_6924; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9997 = 10'h2ff == _dirty_T_1 ? _cache_data_T_6 : _GEN_6925; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9998 = 10'h300 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6926; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_9999 = 10'h301 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6927; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10000 = 10'h302 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6928; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10001 = 10'h303 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6929; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10002 = 10'h304 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6930; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10003 = 10'h305 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6931; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10004 = 10'h306 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6932; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10005 = 10'h307 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6933; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10006 = 10'h308 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6934; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10007 = 10'h309 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6935; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10008 = 10'h30a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6936; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10009 = 10'h30b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6937; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10010 = 10'h30c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6938; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10011 = 10'h30d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6939; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10012 = 10'h30e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6940; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10013 = 10'h30f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6941; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10014 = 10'h310 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6942; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10015 = 10'h311 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6943; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10016 = 10'h312 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6944; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10017 = 10'h313 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6945; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10018 = 10'h314 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6946; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10019 = 10'h315 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6947; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10020 = 10'h316 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6948; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10021 = 10'h317 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6949; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10022 = 10'h318 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6950; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10023 = 10'h319 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6951; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10024 = 10'h31a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6952; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10025 = 10'h31b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6953; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10026 = 10'h31c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6954; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10027 = 10'h31d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6955; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10028 = 10'h31e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6956; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10029 = 10'h31f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6957; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10030 = 10'h320 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6958; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10031 = 10'h321 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6959; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10032 = 10'h322 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6960; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10033 = 10'h323 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6961; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10034 = 10'h324 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6962; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10035 = 10'h325 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6963; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10036 = 10'h326 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6964; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10037 = 10'h327 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6965; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10038 = 10'h328 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6966; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10039 = 10'h329 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6967; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10040 = 10'h32a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6968; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10041 = 10'h32b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6969; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10042 = 10'h32c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6970; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10043 = 10'h32d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6971; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10044 = 10'h32e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6972; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10045 = 10'h32f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6973; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10046 = 10'h330 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6974; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10047 = 10'h331 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6975; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10048 = 10'h332 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6976; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10049 = 10'h333 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6977; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10050 = 10'h334 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6978; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10051 = 10'h335 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6979; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10052 = 10'h336 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6980; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10053 = 10'h337 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6981; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10054 = 10'h338 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6982; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10055 = 10'h339 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6983; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10056 = 10'h33a == _dirty_T_1 ? _cache_data_T_6 : _GEN_6984; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10057 = 10'h33b == _dirty_T_1 ? _cache_data_T_6 : _GEN_6985; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10058 = 10'h33c == _dirty_T_1 ? _cache_data_T_6 : _GEN_6986; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10059 = 10'h33d == _dirty_T_1 ? _cache_data_T_6 : _GEN_6987; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10060 = 10'h33e == _dirty_T_1 ? _cache_data_T_6 : _GEN_6988; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10061 = 10'h33f == _dirty_T_1 ? _cache_data_T_6 : _GEN_6989; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10062 = 10'h340 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6990; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10063 = 10'h341 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6991; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10064 = 10'h342 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6992; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10065 = 10'h343 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6993; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10066 = 10'h344 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6994; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10067 = 10'h345 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6995; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10068 = 10'h346 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6996; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10069 = 10'h347 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6997; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10070 = 10'h348 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6998; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10071 = 10'h349 == _dirty_T_1 ? _cache_data_T_6 : _GEN_6999; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10072 = 10'h34a == _dirty_T_1 ? _cache_data_T_6 : _GEN_7000; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10073 = 10'h34b == _dirty_T_1 ? _cache_data_T_6 : _GEN_7001; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10074 = 10'h34c == _dirty_T_1 ? _cache_data_T_6 : _GEN_7002; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10075 = 10'h34d == _dirty_T_1 ? _cache_data_T_6 : _GEN_7003; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10076 = 10'h34e == _dirty_T_1 ? _cache_data_T_6 : _GEN_7004; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10077 = 10'h34f == _dirty_T_1 ? _cache_data_T_6 : _GEN_7005; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10078 = 10'h350 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7006; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10079 = 10'h351 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7007; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10080 = 10'h352 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7008; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10081 = 10'h353 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7009; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10082 = 10'h354 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7010; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10083 = 10'h355 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7011; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10084 = 10'h356 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7012; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10085 = 10'h357 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7013; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10086 = 10'h358 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7014; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10087 = 10'h359 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7015; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10088 = 10'h35a == _dirty_T_1 ? _cache_data_T_6 : _GEN_7016; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10089 = 10'h35b == _dirty_T_1 ? _cache_data_T_6 : _GEN_7017; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10090 = 10'h35c == _dirty_T_1 ? _cache_data_T_6 : _GEN_7018; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10091 = 10'h35d == _dirty_T_1 ? _cache_data_T_6 : _GEN_7019; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10092 = 10'h35e == _dirty_T_1 ? _cache_data_T_6 : _GEN_7020; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10093 = 10'h35f == _dirty_T_1 ? _cache_data_T_6 : _GEN_7021; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10094 = 10'h360 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7022; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10095 = 10'h361 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7023; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10096 = 10'h362 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7024; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10097 = 10'h363 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7025; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10098 = 10'h364 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7026; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10099 = 10'h365 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7027; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10100 = 10'h366 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7028; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10101 = 10'h367 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7029; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10102 = 10'h368 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7030; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10103 = 10'h369 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7031; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10104 = 10'h36a == _dirty_T_1 ? _cache_data_T_6 : _GEN_7032; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10105 = 10'h36b == _dirty_T_1 ? _cache_data_T_6 : _GEN_7033; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10106 = 10'h36c == _dirty_T_1 ? _cache_data_T_6 : _GEN_7034; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10107 = 10'h36d == _dirty_T_1 ? _cache_data_T_6 : _GEN_7035; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10108 = 10'h36e == _dirty_T_1 ? _cache_data_T_6 : _GEN_7036; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10109 = 10'h36f == _dirty_T_1 ? _cache_data_T_6 : _GEN_7037; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10110 = 10'h370 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7038; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10111 = 10'h371 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7039; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10112 = 10'h372 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7040; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10113 = 10'h373 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7041; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10114 = 10'h374 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7042; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10115 = 10'h375 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7043; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10116 = 10'h376 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7044; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10117 = 10'h377 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7045; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10118 = 10'h378 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7046; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10119 = 10'h379 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7047; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10120 = 10'h37a == _dirty_T_1 ? _cache_data_T_6 : _GEN_7048; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10121 = 10'h37b == _dirty_T_1 ? _cache_data_T_6 : _GEN_7049; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10122 = 10'h37c == _dirty_T_1 ? _cache_data_T_6 : _GEN_7050; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10123 = 10'h37d == _dirty_T_1 ? _cache_data_T_6 : _GEN_7051; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10124 = 10'h37e == _dirty_T_1 ? _cache_data_T_6 : _GEN_7052; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10125 = 10'h37f == _dirty_T_1 ? _cache_data_T_6 : _GEN_7053; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10126 = 10'h380 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7054; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10127 = 10'h381 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7055; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10128 = 10'h382 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7056; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10129 = 10'h383 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7057; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10130 = 10'h384 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7058; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10131 = 10'h385 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7059; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10132 = 10'h386 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7060; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10133 = 10'h387 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7061; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10134 = 10'h388 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7062; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10135 = 10'h389 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7063; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10136 = 10'h38a == _dirty_T_1 ? _cache_data_T_6 : _GEN_7064; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10137 = 10'h38b == _dirty_T_1 ? _cache_data_T_6 : _GEN_7065; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10138 = 10'h38c == _dirty_T_1 ? _cache_data_T_6 : _GEN_7066; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10139 = 10'h38d == _dirty_T_1 ? _cache_data_T_6 : _GEN_7067; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10140 = 10'h38e == _dirty_T_1 ? _cache_data_T_6 : _GEN_7068; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10141 = 10'h38f == _dirty_T_1 ? _cache_data_T_6 : _GEN_7069; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10142 = 10'h390 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7070; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10143 = 10'h391 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7071; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10144 = 10'h392 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7072; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10145 = 10'h393 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7073; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10146 = 10'h394 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7074; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10147 = 10'h395 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7075; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10148 = 10'h396 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7076; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10149 = 10'h397 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7077; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10150 = 10'h398 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7078; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10151 = 10'h399 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7079; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10152 = 10'h39a == _dirty_T_1 ? _cache_data_T_6 : _GEN_7080; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10153 = 10'h39b == _dirty_T_1 ? _cache_data_T_6 : _GEN_7081; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10154 = 10'h39c == _dirty_T_1 ? _cache_data_T_6 : _GEN_7082; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10155 = 10'h39d == _dirty_T_1 ? _cache_data_T_6 : _GEN_7083; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10156 = 10'h39e == _dirty_T_1 ? _cache_data_T_6 : _GEN_7084; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10157 = 10'h39f == _dirty_T_1 ? _cache_data_T_6 : _GEN_7085; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10158 = 10'h3a0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7086; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10159 = 10'h3a1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7087; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10160 = 10'h3a2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7088; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10161 = 10'h3a3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7089; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10162 = 10'h3a4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7090; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10163 = 10'h3a5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7091; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10164 = 10'h3a6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7092; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10165 = 10'h3a7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7093; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10166 = 10'h3a8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7094; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10167 = 10'h3a9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7095; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10168 = 10'h3aa == _dirty_T_1 ? _cache_data_T_6 : _GEN_7096; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10169 = 10'h3ab == _dirty_T_1 ? _cache_data_T_6 : _GEN_7097; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10170 = 10'h3ac == _dirty_T_1 ? _cache_data_T_6 : _GEN_7098; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10171 = 10'h3ad == _dirty_T_1 ? _cache_data_T_6 : _GEN_7099; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10172 = 10'h3ae == _dirty_T_1 ? _cache_data_T_6 : _GEN_7100; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10173 = 10'h3af == _dirty_T_1 ? _cache_data_T_6 : _GEN_7101; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10174 = 10'h3b0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7102; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10175 = 10'h3b1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7103; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10176 = 10'h3b2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7104; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10177 = 10'h3b3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7105; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10178 = 10'h3b4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7106; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10179 = 10'h3b5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7107; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10180 = 10'h3b6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7108; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10181 = 10'h3b7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7109; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10182 = 10'h3b8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7110; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10183 = 10'h3b9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7111; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10184 = 10'h3ba == _dirty_T_1 ? _cache_data_T_6 : _GEN_7112; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10185 = 10'h3bb == _dirty_T_1 ? _cache_data_T_6 : _GEN_7113; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10186 = 10'h3bc == _dirty_T_1 ? _cache_data_T_6 : _GEN_7114; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10187 = 10'h3bd == _dirty_T_1 ? _cache_data_T_6 : _GEN_7115; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10188 = 10'h3be == _dirty_T_1 ? _cache_data_T_6 : _GEN_7116; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10189 = 10'h3bf == _dirty_T_1 ? _cache_data_T_6 : _GEN_7117; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10190 = 10'h3c0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7118; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10191 = 10'h3c1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7119; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10192 = 10'h3c2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7120; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10193 = 10'h3c3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7121; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10194 = 10'h3c4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7122; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10195 = 10'h3c5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7123; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10196 = 10'h3c6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7124; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10197 = 10'h3c7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7125; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10198 = 10'h3c8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7126; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10199 = 10'h3c9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7127; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10200 = 10'h3ca == _dirty_T_1 ? _cache_data_T_6 : _GEN_7128; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10201 = 10'h3cb == _dirty_T_1 ? _cache_data_T_6 : _GEN_7129; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10202 = 10'h3cc == _dirty_T_1 ? _cache_data_T_6 : _GEN_7130; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10203 = 10'h3cd == _dirty_T_1 ? _cache_data_T_6 : _GEN_7131; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10204 = 10'h3ce == _dirty_T_1 ? _cache_data_T_6 : _GEN_7132; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10205 = 10'h3cf == _dirty_T_1 ? _cache_data_T_6 : _GEN_7133; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10206 = 10'h3d0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7134; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10207 = 10'h3d1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7135; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10208 = 10'h3d2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7136; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10209 = 10'h3d3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7137; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10210 = 10'h3d4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7138; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10211 = 10'h3d5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7139; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10212 = 10'h3d6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7140; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10213 = 10'h3d7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7141; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10214 = 10'h3d8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7142; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10215 = 10'h3d9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7143; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10216 = 10'h3da == _dirty_T_1 ? _cache_data_T_6 : _GEN_7144; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10217 = 10'h3db == _dirty_T_1 ? _cache_data_T_6 : _GEN_7145; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10218 = 10'h3dc == _dirty_T_1 ? _cache_data_T_6 : _GEN_7146; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10219 = 10'h3dd == _dirty_T_1 ? _cache_data_T_6 : _GEN_7147; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10220 = 10'h3de == _dirty_T_1 ? _cache_data_T_6 : _GEN_7148; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10221 = 10'h3df == _dirty_T_1 ? _cache_data_T_6 : _GEN_7149; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10222 = 10'h3e0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7150; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10223 = 10'h3e1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7151; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10224 = 10'h3e2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7152; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10225 = 10'h3e3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7153; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10226 = 10'h3e4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7154; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10227 = 10'h3e5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7155; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10228 = 10'h3e6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7156; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10229 = 10'h3e7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7157; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10230 = 10'h3e8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7158; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10231 = 10'h3e9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7159; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10232 = 10'h3ea == _dirty_T_1 ? _cache_data_T_6 : _GEN_7160; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10233 = 10'h3eb == _dirty_T_1 ? _cache_data_T_6 : _GEN_7161; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10234 = 10'h3ec == _dirty_T_1 ? _cache_data_T_6 : _GEN_7162; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10235 = 10'h3ed == _dirty_T_1 ? _cache_data_T_6 : _GEN_7163; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10236 = 10'h3ee == _dirty_T_1 ? _cache_data_T_6 : _GEN_7164; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10237 = 10'h3ef == _dirty_T_1 ? _cache_data_T_6 : _GEN_7165; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10238 = 10'h3f0 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7166; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10239 = 10'h3f1 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7167; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10240 = 10'h3f2 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7168; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10241 = 10'h3f3 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7169; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10242 = 10'h3f4 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7170; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10243 = 10'h3f5 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7171; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10244 = 10'h3f6 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7172; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10245 = 10'h3f7 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7173; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10246 = 10'h3f8 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7174; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10247 = 10'h3f9 == _dirty_T_1 ? _cache_data_T_6 : _GEN_7175; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10248 = 10'h3fa == _dirty_T_1 ? _cache_data_T_6 : _GEN_7176; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10249 = 10'h3fb == _dirty_T_1 ? _cache_data_T_6 : _GEN_7177; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10250 = 10'h3fc == _dirty_T_1 ? _cache_data_T_6 : _GEN_7178; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10251 = 10'h3fd == _dirty_T_1 ? _cache_data_T_6 : _GEN_7179; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10252 = 10'h3fe == _dirty_T_1 ? _cache_data_T_6 : _GEN_7180; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10253 = 10'h3ff == _dirty_T_1 ? _cache_data_T_6 : _GEN_7181; // @[icache.scala 136:{33,33}]
  wire [184:0] _GEN_10254 = replace & io_inst_sram_data_ok ? _GEN_9230 : _GEN_6158; // @[icache.scala 135:42]
  wire [184:0] _GEN_10255 = replace & io_inst_sram_data_ok ? _GEN_9231 : _GEN_6159; // @[icache.scala 135:42]
  wire [184:0] _GEN_10256 = replace & io_inst_sram_data_ok ? _GEN_9232 : _GEN_6160; // @[icache.scala 135:42]
  wire [184:0] _GEN_10257 = replace & io_inst_sram_data_ok ? _GEN_9233 : _GEN_6161; // @[icache.scala 135:42]
  wire [184:0] _GEN_10258 = replace & io_inst_sram_data_ok ? _GEN_9234 : _GEN_6162; // @[icache.scala 135:42]
  wire [184:0] _GEN_10259 = replace & io_inst_sram_data_ok ? _GEN_9235 : _GEN_6163; // @[icache.scala 135:42]
  wire [184:0] _GEN_10260 = replace & io_inst_sram_data_ok ? _GEN_9236 : _GEN_6164; // @[icache.scala 135:42]
  wire [184:0] _GEN_10261 = replace & io_inst_sram_data_ok ? _GEN_9237 : _GEN_6165; // @[icache.scala 135:42]
  wire [184:0] _GEN_10262 = replace & io_inst_sram_data_ok ? _GEN_9238 : _GEN_6166; // @[icache.scala 135:42]
  wire [184:0] _GEN_10263 = replace & io_inst_sram_data_ok ? _GEN_9239 : _GEN_6167; // @[icache.scala 135:42]
  wire [184:0] _GEN_10264 = replace & io_inst_sram_data_ok ? _GEN_9240 : _GEN_6168; // @[icache.scala 135:42]
  wire [184:0] _GEN_10265 = replace & io_inst_sram_data_ok ? _GEN_9241 : _GEN_6169; // @[icache.scala 135:42]
  wire [184:0] _GEN_10266 = replace & io_inst_sram_data_ok ? _GEN_9242 : _GEN_6170; // @[icache.scala 135:42]
  wire [184:0] _GEN_10267 = replace & io_inst_sram_data_ok ? _GEN_9243 : _GEN_6171; // @[icache.scala 135:42]
  wire [184:0] _GEN_10268 = replace & io_inst_sram_data_ok ? _GEN_9244 : _GEN_6172; // @[icache.scala 135:42]
  wire [184:0] _GEN_10269 = replace & io_inst_sram_data_ok ? _GEN_9245 : _GEN_6173; // @[icache.scala 135:42]
  wire [184:0] _GEN_10270 = replace & io_inst_sram_data_ok ? _GEN_9246 : _GEN_6174; // @[icache.scala 135:42]
  wire [184:0] _GEN_10271 = replace & io_inst_sram_data_ok ? _GEN_9247 : _GEN_6175; // @[icache.scala 135:42]
  wire [184:0] _GEN_10272 = replace & io_inst_sram_data_ok ? _GEN_9248 : _GEN_6176; // @[icache.scala 135:42]
  wire [184:0] _GEN_10273 = replace & io_inst_sram_data_ok ? _GEN_9249 : _GEN_6177; // @[icache.scala 135:42]
  wire [184:0] _GEN_10274 = replace & io_inst_sram_data_ok ? _GEN_9250 : _GEN_6178; // @[icache.scala 135:42]
  wire [184:0] _GEN_10275 = replace & io_inst_sram_data_ok ? _GEN_9251 : _GEN_6179; // @[icache.scala 135:42]
  wire [184:0] _GEN_10276 = replace & io_inst_sram_data_ok ? _GEN_9252 : _GEN_6180; // @[icache.scala 135:42]
  wire [184:0] _GEN_10277 = replace & io_inst_sram_data_ok ? _GEN_9253 : _GEN_6181; // @[icache.scala 135:42]
  wire [184:0] _GEN_10278 = replace & io_inst_sram_data_ok ? _GEN_9254 : _GEN_6182; // @[icache.scala 135:42]
  wire [184:0] _GEN_10279 = replace & io_inst_sram_data_ok ? _GEN_9255 : _GEN_6183; // @[icache.scala 135:42]
  wire [184:0] _GEN_10280 = replace & io_inst_sram_data_ok ? _GEN_9256 : _GEN_6184; // @[icache.scala 135:42]
  wire [184:0] _GEN_10281 = replace & io_inst_sram_data_ok ? _GEN_9257 : _GEN_6185; // @[icache.scala 135:42]
  wire [184:0] _GEN_10282 = replace & io_inst_sram_data_ok ? _GEN_9258 : _GEN_6186; // @[icache.scala 135:42]
  wire [184:0] _GEN_10283 = replace & io_inst_sram_data_ok ? _GEN_9259 : _GEN_6187; // @[icache.scala 135:42]
  wire [184:0] _GEN_10284 = replace & io_inst_sram_data_ok ? _GEN_9260 : _GEN_6188; // @[icache.scala 135:42]
  wire [184:0] _GEN_10285 = replace & io_inst_sram_data_ok ? _GEN_9261 : _GEN_6189; // @[icache.scala 135:42]
  wire [184:0] _GEN_10286 = replace & io_inst_sram_data_ok ? _GEN_9262 : _GEN_6190; // @[icache.scala 135:42]
  wire [184:0] _GEN_10287 = replace & io_inst_sram_data_ok ? _GEN_9263 : _GEN_6191; // @[icache.scala 135:42]
  wire [184:0] _GEN_10288 = replace & io_inst_sram_data_ok ? _GEN_9264 : _GEN_6192; // @[icache.scala 135:42]
  wire [184:0] _GEN_10289 = replace & io_inst_sram_data_ok ? _GEN_9265 : _GEN_6193; // @[icache.scala 135:42]
  wire [184:0] _GEN_10290 = replace & io_inst_sram_data_ok ? _GEN_9266 : _GEN_6194; // @[icache.scala 135:42]
  wire [184:0] _GEN_10291 = replace & io_inst_sram_data_ok ? _GEN_9267 : _GEN_6195; // @[icache.scala 135:42]
  wire [184:0] _GEN_10292 = replace & io_inst_sram_data_ok ? _GEN_9268 : _GEN_6196; // @[icache.scala 135:42]
  wire [184:0] _GEN_10293 = replace & io_inst_sram_data_ok ? _GEN_9269 : _GEN_6197; // @[icache.scala 135:42]
  wire [184:0] _GEN_10294 = replace & io_inst_sram_data_ok ? _GEN_9270 : _GEN_6198; // @[icache.scala 135:42]
  wire [184:0] _GEN_10295 = replace & io_inst_sram_data_ok ? _GEN_9271 : _GEN_6199; // @[icache.scala 135:42]
  wire [184:0] _GEN_10296 = replace & io_inst_sram_data_ok ? _GEN_9272 : _GEN_6200; // @[icache.scala 135:42]
  wire [184:0] _GEN_10297 = replace & io_inst_sram_data_ok ? _GEN_9273 : _GEN_6201; // @[icache.scala 135:42]
  wire [184:0] _GEN_10298 = replace & io_inst_sram_data_ok ? _GEN_9274 : _GEN_6202; // @[icache.scala 135:42]
  wire [184:0] _GEN_10299 = replace & io_inst_sram_data_ok ? _GEN_9275 : _GEN_6203; // @[icache.scala 135:42]
  wire [184:0] _GEN_10300 = replace & io_inst_sram_data_ok ? _GEN_9276 : _GEN_6204; // @[icache.scala 135:42]
  wire [184:0] _GEN_10301 = replace & io_inst_sram_data_ok ? _GEN_9277 : _GEN_6205; // @[icache.scala 135:42]
  wire [184:0] _GEN_10302 = replace & io_inst_sram_data_ok ? _GEN_9278 : _GEN_6206; // @[icache.scala 135:42]
  wire [184:0] _GEN_10303 = replace & io_inst_sram_data_ok ? _GEN_9279 : _GEN_6207; // @[icache.scala 135:42]
  wire [184:0] _GEN_10304 = replace & io_inst_sram_data_ok ? _GEN_9280 : _GEN_6208; // @[icache.scala 135:42]
  wire [184:0] _GEN_10305 = replace & io_inst_sram_data_ok ? _GEN_9281 : _GEN_6209; // @[icache.scala 135:42]
  wire [184:0] _GEN_10306 = replace & io_inst_sram_data_ok ? _GEN_9282 : _GEN_6210; // @[icache.scala 135:42]
  wire [184:0] _GEN_10307 = replace & io_inst_sram_data_ok ? _GEN_9283 : _GEN_6211; // @[icache.scala 135:42]
  wire [184:0] _GEN_10308 = replace & io_inst_sram_data_ok ? _GEN_9284 : _GEN_6212; // @[icache.scala 135:42]
  wire [184:0] _GEN_10309 = replace & io_inst_sram_data_ok ? _GEN_9285 : _GEN_6213; // @[icache.scala 135:42]
  wire [184:0] _GEN_10310 = replace & io_inst_sram_data_ok ? _GEN_9286 : _GEN_6214; // @[icache.scala 135:42]
  wire [184:0] _GEN_10311 = replace & io_inst_sram_data_ok ? _GEN_9287 : _GEN_6215; // @[icache.scala 135:42]
  wire [184:0] _GEN_10312 = replace & io_inst_sram_data_ok ? _GEN_9288 : _GEN_6216; // @[icache.scala 135:42]
  wire [184:0] _GEN_10313 = replace & io_inst_sram_data_ok ? _GEN_9289 : _GEN_6217; // @[icache.scala 135:42]
  wire [184:0] _GEN_10314 = replace & io_inst_sram_data_ok ? _GEN_9290 : _GEN_6218; // @[icache.scala 135:42]
  wire [184:0] _GEN_10315 = replace & io_inst_sram_data_ok ? _GEN_9291 : _GEN_6219; // @[icache.scala 135:42]
  wire [184:0] _GEN_10316 = replace & io_inst_sram_data_ok ? _GEN_9292 : _GEN_6220; // @[icache.scala 135:42]
  wire [184:0] _GEN_10317 = replace & io_inst_sram_data_ok ? _GEN_9293 : _GEN_6221; // @[icache.scala 135:42]
  wire [184:0] _GEN_10318 = replace & io_inst_sram_data_ok ? _GEN_9294 : _GEN_6222; // @[icache.scala 135:42]
  wire [184:0] _GEN_10319 = replace & io_inst_sram_data_ok ? _GEN_9295 : _GEN_6223; // @[icache.scala 135:42]
  wire [184:0] _GEN_10320 = replace & io_inst_sram_data_ok ? _GEN_9296 : _GEN_6224; // @[icache.scala 135:42]
  wire [184:0] _GEN_10321 = replace & io_inst_sram_data_ok ? _GEN_9297 : _GEN_6225; // @[icache.scala 135:42]
  wire [184:0] _GEN_10322 = replace & io_inst_sram_data_ok ? _GEN_9298 : _GEN_6226; // @[icache.scala 135:42]
  wire [184:0] _GEN_10323 = replace & io_inst_sram_data_ok ? _GEN_9299 : _GEN_6227; // @[icache.scala 135:42]
  wire [184:0] _GEN_10324 = replace & io_inst_sram_data_ok ? _GEN_9300 : _GEN_6228; // @[icache.scala 135:42]
  wire [184:0] _GEN_10325 = replace & io_inst_sram_data_ok ? _GEN_9301 : _GEN_6229; // @[icache.scala 135:42]
  wire [184:0] _GEN_10326 = replace & io_inst_sram_data_ok ? _GEN_9302 : _GEN_6230; // @[icache.scala 135:42]
  wire [184:0] _GEN_10327 = replace & io_inst_sram_data_ok ? _GEN_9303 : _GEN_6231; // @[icache.scala 135:42]
  wire [184:0] _GEN_10328 = replace & io_inst_sram_data_ok ? _GEN_9304 : _GEN_6232; // @[icache.scala 135:42]
  wire [184:0] _GEN_10329 = replace & io_inst_sram_data_ok ? _GEN_9305 : _GEN_6233; // @[icache.scala 135:42]
  wire [184:0] _GEN_10330 = replace & io_inst_sram_data_ok ? _GEN_9306 : _GEN_6234; // @[icache.scala 135:42]
  wire [184:0] _GEN_10331 = replace & io_inst_sram_data_ok ? _GEN_9307 : _GEN_6235; // @[icache.scala 135:42]
  wire [184:0] _GEN_10332 = replace & io_inst_sram_data_ok ? _GEN_9308 : _GEN_6236; // @[icache.scala 135:42]
  wire [184:0] _GEN_10333 = replace & io_inst_sram_data_ok ? _GEN_9309 : _GEN_6237; // @[icache.scala 135:42]
  wire [184:0] _GEN_10334 = replace & io_inst_sram_data_ok ? _GEN_9310 : _GEN_6238; // @[icache.scala 135:42]
  wire [184:0] _GEN_10335 = replace & io_inst_sram_data_ok ? _GEN_9311 : _GEN_6239; // @[icache.scala 135:42]
  wire [184:0] _GEN_10336 = replace & io_inst_sram_data_ok ? _GEN_9312 : _GEN_6240; // @[icache.scala 135:42]
  wire [184:0] _GEN_10337 = replace & io_inst_sram_data_ok ? _GEN_9313 : _GEN_6241; // @[icache.scala 135:42]
  wire [184:0] _GEN_10338 = replace & io_inst_sram_data_ok ? _GEN_9314 : _GEN_6242; // @[icache.scala 135:42]
  wire [184:0] _GEN_10339 = replace & io_inst_sram_data_ok ? _GEN_9315 : _GEN_6243; // @[icache.scala 135:42]
  wire [184:0] _GEN_10340 = replace & io_inst_sram_data_ok ? _GEN_9316 : _GEN_6244; // @[icache.scala 135:42]
  wire [184:0] _GEN_10341 = replace & io_inst_sram_data_ok ? _GEN_9317 : _GEN_6245; // @[icache.scala 135:42]
  wire [184:0] _GEN_10342 = replace & io_inst_sram_data_ok ? _GEN_9318 : _GEN_6246; // @[icache.scala 135:42]
  wire [184:0] _GEN_10343 = replace & io_inst_sram_data_ok ? _GEN_9319 : _GEN_6247; // @[icache.scala 135:42]
  wire [184:0] _GEN_10344 = replace & io_inst_sram_data_ok ? _GEN_9320 : _GEN_6248; // @[icache.scala 135:42]
  wire [184:0] _GEN_10345 = replace & io_inst_sram_data_ok ? _GEN_9321 : _GEN_6249; // @[icache.scala 135:42]
  wire [184:0] _GEN_10346 = replace & io_inst_sram_data_ok ? _GEN_9322 : _GEN_6250; // @[icache.scala 135:42]
  wire [184:0] _GEN_10347 = replace & io_inst_sram_data_ok ? _GEN_9323 : _GEN_6251; // @[icache.scala 135:42]
  wire [184:0] _GEN_10348 = replace & io_inst_sram_data_ok ? _GEN_9324 : _GEN_6252; // @[icache.scala 135:42]
  wire [184:0] _GEN_10349 = replace & io_inst_sram_data_ok ? _GEN_9325 : _GEN_6253; // @[icache.scala 135:42]
  wire [184:0] _GEN_10350 = replace & io_inst_sram_data_ok ? _GEN_9326 : _GEN_6254; // @[icache.scala 135:42]
  wire [184:0] _GEN_10351 = replace & io_inst_sram_data_ok ? _GEN_9327 : _GEN_6255; // @[icache.scala 135:42]
  wire [184:0] _GEN_10352 = replace & io_inst_sram_data_ok ? _GEN_9328 : _GEN_6256; // @[icache.scala 135:42]
  wire [184:0] _GEN_10353 = replace & io_inst_sram_data_ok ? _GEN_9329 : _GEN_6257; // @[icache.scala 135:42]
  wire [184:0] _GEN_10354 = replace & io_inst_sram_data_ok ? _GEN_9330 : _GEN_6258; // @[icache.scala 135:42]
  wire [184:0] _GEN_10355 = replace & io_inst_sram_data_ok ? _GEN_9331 : _GEN_6259; // @[icache.scala 135:42]
  wire [184:0] _GEN_10356 = replace & io_inst_sram_data_ok ? _GEN_9332 : _GEN_6260; // @[icache.scala 135:42]
  wire [184:0] _GEN_10357 = replace & io_inst_sram_data_ok ? _GEN_9333 : _GEN_6261; // @[icache.scala 135:42]
  wire [184:0] _GEN_10358 = replace & io_inst_sram_data_ok ? _GEN_9334 : _GEN_6262; // @[icache.scala 135:42]
  wire [184:0] _GEN_10359 = replace & io_inst_sram_data_ok ? _GEN_9335 : _GEN_6263; // @[icache.scala 135:42]
  wire [184:0] _GEN_10360 = replace & io_inst_sram_data_ok ? _GEN_9336 : _GEN_6264; // @[icache.scala 135:42]
  wire [184:0] _GEN_10361 = replace & io_inst_sram_data_ok ? _GEN_9337 : _GEN_6265; // @[icache.scala 135:42]
  wire [184:0] _GEN_10362 = replace & io_inst_sram_data_ok ? _GEN_9338 : _GEN_6266; // @[icache.scala 135:42]
  wire [184:0] _GEN_10363 = replace & io_inst_sram_data_ok ? _GEN_9339 : _GEN_6267; // @[icache.scala 135:42]
  wire [184:0] _GEN_10364 = replace & io_inst_sram_data_ok ? _GEN_9340 : _GEN_6268; // @[icache.scala 135:42]
  wire [184:0] _GEN_10365 = replace & io_inst_sram_data_ok ? _GEN_9341 : _GEN_6269; // @[icache.scala 135:42]
  wire [184:0] _GEN_10366 = replace & io_inst_sram_data_ok ? _GEN_9342 : _GEN_6270; // @[icache.scala 135:42]
  wire [184:0] _GEN_10367 = replace & io_inst_sram_data_ok ? _GEN_9343 : _GEN_6271; // @[icache.scala 135:42]
  wire [184:0] _GEN_10368 = replace & io_inst_sram_data_ok ? _GEN_9344 : _GEN_6272; // @[icache.scala 135:42]
  wire [184:0] _GEN_10369 = replace & io_inst_sram_data_ok ? _GEN_9345 : _GEN_6273; // @[icache.scala 135:42]
  wire [184:0] _GEN_10370 = replace & io_inst_sram_data_ok ? _GEN_9346 : _GEN_6274; // @[icache.scala 135:42]
  wire [184:0] _GEN_10371 = replace & io_inst_sram_data_ok ? _GEN_9347 : _GEN_6275; // @[icache.scala 135:42]
  wire [184:0] _GEN_10372 = replace & io_inst_sram_data_ok ? _GEN_9348 : _GEN_6276; // @[icache.scala 135:42]
  wire [184:0] _GEN_10373 = replace & io_inst_sram_data_ok ? _GEN_9349 : _GEN_6277; // @[icache.scala 135:42]
  wire [184:0] _GEN_10374 = replace & io_inst_sram_data_ok ? _GEN_9350 : _GEN_6278; // @[icache.scala 135:42]
  wire [184:0] _GEN_10375 = replace & io_inst_sram_data_ok ? _GEN_9351 : _GEN_6279; // @[icache.scala 135:42]
  wire [184:0] _GEN_10376 = replace & io_inst_sram_data_ok ? _GEN_9352 : _GEN_6280; // @[icache.scala 135:42]
  wire [184:0] _GEN_10377 = replace & io_inst_sram_data_ok ? _GEN_9353 : _GEN_6281; // @[icache.scala 135:42]
  wire [184:0] _GEN_10378 = replace & io_inst_sram_data_ok ? _GEN_9354 : _GEN_6282; // @[icache.scala 135:42]
  wire [184:0] _GEN_10379 = replace & io_inst_sram_data_ok ? _GEN_9355 : _GEN_6283; // @[icache.scala 135:42]
  wire [184:0] _GEN_10380 = replace & io_inst_sram_data_ok ? _GEN_9356 : _GEN_6284; // @[icache.scala 135:42]
  wire [184:0] _GEN_10381 = replace & io_inst_sram_data_ok ? _GEN_9357 : _GEN_6285; // @[icache.scala 135:42]
  wire [184:0] _GEN_10382 = replace & io_inst_sram_data_ok ? _GEN_9358 : _GEN_6286; // @[icache.scala 135:42]
  wire [184:0] _GEN_10383 = replace & io_inst_sram_data_ok ? _GEN_9359 : _GEN_6287; // @[icache.scala 135:42]
  wire [184:0] _GEN_10384 = replace & io_inst_sram_data_ok ? _GEN_9360 : _GEN_6288; // @[icache.scala 135:42]
  wire [184:0] _GEN_10385 = replace & io_inst_sram_data_ok ? _GEN_9361 : _GEN_6289; // @[icache.scala 135:42]
  wire [184:0] _GEN_10386 = replace & io_inst_sram_data_ok ? _GEN_9362 : _GEN_6290; // @[icache.scala 135:42]
  wire [184:0] _GEN_10387 = replace & io_inst_sram_data_ok ? _GEN_9363 : _GEN_6291; // @[icache.scala 135:42]
  wire [184:0] _GEN_10388 = replace & io_inst_sram_data_ok ? _GEN_9364 : _GEN_6292; // @[icache.scala 135:42]
  wire [184:0] _GEN_10389 = replace & io_inst_sram_data_ok ? _GEN_9365 : _GEN_6293; // @[icache.scala 135:42]
  wire [184:0] _GEN_10390 = replace & io_inst_sram_data_ok ? _GEN_9366 : _GEN_6294; // @[icache.scala 135:42]
  wire [184:0] _GEN_10391 = replace & io_inst_sram_data_ok ? _GEN_9367 : _GEN_6295; // @[icache.scala 135:42]
  wire [184:0] _GEN_10392 = replace & io_inst_sram_data_ok ? _GEN_9368 : _GEN_6296; // @[icache.scala 135:42]
  wire [184:0] _GEN_10393 = replace & io_inst_sram_data_ok ? _GEN_9369 : _GEN_6297; // @[icache.scala 135:42]
  wire [184:0] _GEN_10394 = replace & io_inst_sram_data_ok ? _GEN_9370 : _GEN_6298; // @[icache.scala 135:42]
  wire [184:0] _GEN_10395 = replace & io_inst_sram_data_ok ? _GEN_9371 : _GEN_6299; // @[icache.scala 135:42]
  wire [184:0] _GEN_10396 = replace & io_inst_sram_data_ok ? _GEN_9372 : _GEN_6300; // @[icache.scala 135:42]
  wire [184:0] _GEN_10397 = replace & io_inst_sram_data_ok ? _GEN_9373 : _GEN_6301; // @[icache.scala 135:42]
  wire [184:0] _GEN_10398 = replace & io_inst_sram_data_ok ? _GEN_9374 : _GEN_6302; // @[icache.scala 135:42]
  wire [184:0] _GEN_10399 = replace & io_inst_sram_data_ok ? _GEN_9375 : _GEN_6303; // @[icache.scala 135:42]
  wire [184:0] _GEN_10400 = replace & io_inst_sram_data_ok ? _GEN_9376 : _GEN_6304; // @[icache.scala 135:42]
  wire [184:0] _GEN_10401 = replace & io_inst_sram_data_ok ? _GEN_9377 : _GEN_6305; // @[icache.scala 135:42]
  wire [184:0] _GEN_10402 = replace & io_inst_sram_data_ok ? _GEN_9378 : _GEN_6306; // @[icache.scala 135:42]
  wire [184:0] _GEN_10403 = replace & io_inst_sram_data_ok ? _GEN_9379 : _GEN_6307; // @[icache.scala 135:42]
  wire [184:0] _GEN_10404 = replace & io_inst_sram_data_ok ? _GEN_9380 : _GEN_6308; // @[icache.scala 135:42]
  wire [184:0] _GEN_10405 = replace & io_inst_sram_data_ok ? _GEN_9381 : _GEN_6309; // @[icache.scala 135:42]
  wire [184:0] _GEN_10406 = replace & io_inst_sram_data_ok ? _GEN_9382 : _GEN_6310; // @[icache.scala 135:42]
  wire [184:0] _GEN_10407 = replace & io_inst_sram_data_ok ? _GEN_9383 : _GEN_6311; // @[icache.scala 135:42]
  wire [184:0] _GEN_10408 = replace & io_inst_sram_data_ok ? _GEN_9384 : _GEN_6312; // @[icache.scala 135:42]
  wire [184:0] _GEN_10409 = replace & io_inst_sram_data_ok ? _GEN_9385 : _GEN_6313; // @[icache.scala 135:42]
  wire [184:0] _GEN_10410 = replace & io_inst_sram_data_ok ? _GEN_9386 : _GEN_6314; // @[icache.scala 135:42]
  wire [184:0] _GEN_10411 = replace & io_inst_sram_data_ok ? _GEN_9387 : _GEN_6315; // @[icache.scala 135:42]
  wire [184:0] _GEN_10412 = replace & io_inst_sram_data_ok ? _GEN_9388 : _GEN_6316; // @[icache.scala 135:42]
  wire [184:0] _GEN_10413 = replace & io_inst_sram_data_ok ? _GEN_9389 : _GEN_6317; // @[icache.scala 135:42]
  wire [184:0] _GEN_10414 = replace & io_inst_sram_data_ok ? _GEN_9390 : _GEN_6318; // @[icache.scala 135:42]
  wire [184:0] _GEN_10415 = replace & io_inst_sram_data_ok ? _GEN_9391 : _GEN_6319; // @[icache.scala 135:42]
  wire [184:0] _GEN_10416 = replace & io_inst_sram_data_ok ? _GEN_9392 : _GEN_6320; // @[icache.scala 135:42]
  wire [184:0] _GEN_10417 = replace & io_inst_sram_data_ok ? _GEN_9393 : _GEN_6321; // @[icache.scala 135:42]
  wire [184:0] _GEN_10418 = replace & io_inst_sram_data_ok ? _GEN_9394 : _GEN_6322; // @[icache.scala 135:42]
  wire [184:0] _GEN_10419 = replace & io_inst_sram_data_ok ? _GEN_9395 : _GEN_6323; // @[icache.scala 135:42]
  wire [184:0] _GEN_10420 = replace & io_inst_sram_data_ok ? _GEN_9396 : _GEN_6324; // @[icache.scala 135:42]
  wire [184:0] _GEN_10421 = replace & io_inst_sram_data_ok ? _GEN_9397 : _GEN_6325; // @[icache.scala 135:42]
  wire [184:0] _GEN_10422 = replace & io_inst_sram_data_ok ? _GEN_9398 : _GEN_6326; // @[icache.scala 135:42]
  wire [184:0] _GEN_10423 = replace & io_inst_sram_data_ok ? _GEN_9399 : _GEN_6327; // @[icache.scala 135:42]
  wire [184:0] _GEN_10424 = replace & io_inst_sram_data_ok ? _GEN_9400 : _GEN_6328; // @[icache.scala 135:42]
  wire [184:0] _GEN_10425 = replace & io_inst_sram_data_ok ? _GEN_9401 : _GEN_6329; // @[icache.scala 135:42]
  wire [184:0] _GEN_10426 = replace & io_inst_sram_data_ok ? _GEN_9402 : _GEN_6330; // @[icache.scala 135:42]
  wire [184:0] _GEN_10427 = replace & io_inst_sram_data_ok ? _GEN_9403 : _GEN_6331; // @[icache.scala 135:42]
  wire [184:0] _GEN_10428 = replace & io_inst_sram_data_ok ? _GEN_9404 : _GEN_6332; // @[icache.scala 135:42]
  wire [184:0] _GEN_10429 = replace & io_inst_sram_data_ok ? _GEN_9405 : _GEN_6333; // @[icache.scala 135:42]
  wire [184:0] _GEN_10430 = replace & io_inst_sram_data_ok ? _GEN_9406 : _GEN_6334; // @[icache.scala 135:42]
  wire [184:0] _GEN_10431 = replace & io_inst_sram_data_ok ? _GEN_9407 : _GEN_6335; // @[icache.scala 135:42]
  wire [184:0] _GEN_10432 = replace & io_inst_sram_data_ok ? _GEN_9408 : _GEN_6336; // @[icache.scala 135:42]
  wire [184:0] _GEN_10433 = replace & io_inst_sram_data_ok ? _GEN_9409 : _GEN_6337; // @[icache.scala 135:42]
  wire [184:0] _GEN_10434 = replace & io_inst_sram_data_ok ? _GEN_9410 : _GEN_6338; // @[icache.scala 135:42]
  wire [184:0] _GEN_10435 = replace & io_inst_sram_data_ok ? _GEN_9411 : _GEN_6339; // @[icache.scala 135:42]
  wire [184:0] _GEN_10436 = replace & io_inst_sram_data_ok ? _GEN_9412 : _GEN_6340; // @[icache.scala 135:42]
  wire [184:0] _GEN_10437 = replace & io_inst_sram_data_ok ? _GEN_9413 : _GEN_6341; // @[icache.scala 135:42]
  wire [184:0] _GEN_10438 = replace & io_inst_sram_data_ok ? _GEN_9414 : _GEN_6342; // @[icache.scala 135:42]
  wire [184:0] _GEN_10439 = replace & io_inst_sram_data_ok ? _GEN_9415 : _GEN_6343; // @[icache.scala 135:42]
  wire [184:0] _GEN_10440 = replace & io_inst_sram_data_ok ? _GEN_9416 : _GEN_6344; // @[icache.scala 135:42]
  wire [184:0] _GEN_10441 = replace & io_inst_sram_data_ok ? _GEN_9417 : _GEN_6345; // @[icache.scala 135:42]
  wire [184:0] _GEN_10442 = replace & io_inst_sram_data_ok ? _GEN_9418 : _GEN_6346; // @[icache.scala 135:42]
  wire [184:0] _GEN_10443 = replace & io_inst_sram_data_ok ? _GEN_9419 : _GEN_6347; // @[icache.scala 135:42]
  wire [184:0] _GEN_10444 = replace & io_inst_sram_data_ok ? _GEN_9420 : _GEN_6348; // @[icache.scala 135:42]
  wire [184:0] _GEN_10445 = replace & io_inst_sram_data_ok ? _GEN_9421 : _GEN_6349; // @[icache.scala 135:42]
  wire [184:0] _GEN_10446 = replace & io_inst_sram_data_ok ? _GEN_9422 : _GEN_6350; // @[icache.scala 135:42]
  wire [184:0] _GEN_10447 = replace & io_inst_sram_data_ok ? _GEN_9423 : _GEN_6351; // @[icache.scala 135:42]
  wire [184:0] _GEN_10448 = replace & io_inst_sram_data_ok ? _GEN_9424 : _GEN_6352; // @[icache.scala 135:42]
  wire [184:0] _GEN_10449 = replace & io_inst_sram_data_ok ? _GEN_9425 : _GEN_6353; // @[icache.scala 135:42]
  wire [184:0] _GEN_10450 = replace & io_inst_sram_data_ok ? _GEN_9426 : _GEN_6354; // @[icache.scala 135:42]
  wire [184:0] _GEN_10451 = replace & io_inst_sram_data_ok ? _GEN_9427 : _GEN_6355; // @[icache.scala 135:42]
  wire [184:0] _GEN_10452 = replace & io_inst_sram_data_ok ? _GEN_9428 : _GEN_6356; // @[icache.scala 135:42]
  wire [184:0] _GEN_10453 = replace & io_inst_sram_data_ok ? _GEN_9429 : _GEN_6357; // @[icache.scala 135:42]
  wire [184:0] _GEN_10454 = replace & io_inst_sram_data_ok ? _GEN_9430 : _GEN_6358; // @[icache.scala 135:42]
  wire [184:0] _GEN_10455 = replace & io_inst_sram_data_ok ? _GEN_9431 : _GEN_6359; // @[icache.scala 135:42]
  wire [184:0] _GEN_10456 = replace & io_inst_sram_data_ok ? _GEN_9432 : _GEN_6360; // @[icache.scala 135:42]
  wire [184:0] _GEN_10457 = replace & io_inst_sram_data_ok ? _GEN_9433 : _GEN_6361; // @[icache.scala 135:42]
  wire [184:0] _GEN_10458 = replace & io_inst_sram_data_ok ? _GEN_9434 : _GEN_6362; // @[icache.scala 135:42]
  wire [184:0] _GEN_10459 = replace & io_inst_sram_data_ok ? _GEN_9435 : _GEN_6363; // @[icache.scala 135:42]
  wire [184:0] _GEN_10460 = replace & io_inst_sram_data_ok ? _GEN_9436 : _GEN_6364; // @[icache.scala 135:42]
  wire [184:0] _GEN_10461 = replace & io_inst_sram_data_ok ? _GEN_9437 : _GEN_6365; // @[icache.scala 135:42]
  wire [184:0] _GEN_10462 = replace & io_inst_sram_data_ok ? _GEN_9438 : _GEN_6366; // @[icache.scala 135:42]
  wire [184:0] _GEN_10463 = replace & io_inst_sram_data_ok ? _GEN_9439 : _GEN_6367; // @[icache.scala 135:42]
  wire [184:0] _GEN_10464 = replace & io_inst_sram_data_ok ? _GEN_9440 : _GEN_6368; // @[icache.scala 135:42]
  wire [184:0] _GEN_10465 = replace & io_inst_sram_data_ok ? _GEN_9441 : _GEN_6369; // @[icache.scala 135:42]
  wire [184:0] _GEN_10466 = replace & io_inst_sram_data_ok ? _GEN_9442 : _GEN_6370; // @[icache.scala 135:42]
  wire [184:0] _GEN_10467 = replace & io_inst_sram_data_ok ? _GEN_9443 : _GEN_6371; // @[icache.scala 135:42]
  wire [184:0] _GEN_10468 = replace & io_inst_sram_data_ok ? _GEN_9444 : _GEN_6372; // @[icache.scala 135:42]
  wire [184:0] _GEN_10469 = replace & io_inst_sram_data_ok ? _GEN_9445 : _GEN_6373; // @[icache.scala 135:42]
  wire [184:0] _GEN_10470 = replace & io_inst_sram_data_ok ? _GEN_9446 : _GEN_6374; // @[icache.scala 135:42]
  wire [184:0] _GEN_10471 = replace & io_inst_sram_data_ok ? _GEN_9447 : _GEN_6375; // @[icache.scala 135:42]
  wire [184:0] _GEN_10472 = replace & io_inst_sram_data_ok ? _GEN_9448 : _GEN_6376; // @[icache.scala 135:42]
  wire [184:0] _GEN_10473 = replace & io_inst_sram_data_ok ? _GEN_9449 : _GEN_6377; // @[icache.scala 135:42]
  wire [184:0] _GEN_10474 = replace & io_inst_sram_data_ok ? _GEN_9450 : _GEN_6378; // @[icache.scala 135:42]
  wire [184:0] _GEN_10475 = replace & io_inst_sram_data_ok ? _GEN_9451 : _GEN_6379; // @[icache.scala 135:42]
  wire [184:0] _GEN_10476 = replace & io_inst_sram_data_ok ? _GEN_9452 : _GEN_6380; // @[icache.scala 135:42]
  wire [184:0] _GEN_10477 = replace & io_inst_sram_data_ok ? _GEN_9453 : _GEN_6381; // @[icache.scala 135:42]
  wire [184:0] _GEN_10478 = replace & io_inst_sram_data_ok ? _GEN_9454 : _GEN_6382; // @[icache.scala 135:42]
  wire [184:0] _GEN_10479 = replace & io_inst_sram_data_ok ? _GEN_9455 : _GEN_6383; // @[icache.scala 135:42]
  wire [184:0] _GEN_10480 = replace & io_inst_sram_data_ok ? _GEN_9456 : _GEN_6384; // @[icache.scala 135:42]
  wire [184:0] _GEN_10481 = replace & io_inst_sram_data_ok ? _GEN_9457 : _GEN_6385; // @[icache.scala 135:42]
  wire [184:0] _GEN_10482 = replace & io_inst_sram_data_ok ? _GEN_9458 : _GEN_6386; // @[icache.scala 135:42]
  wire [184:0] _GEN_10483 = replace & io_inst_sram_data_ok ? _GEN_9459 : _GEN_6387; // @[icache.scala 135:42]
  wire [184:0] _GEN_10484 = replace & io_inst_sram_data_ok ? _GEN_9460 : _GEN_6388; // @[icache.scala 135:42]
  wire [184:0] _GEN_10485 = replace & io_inst_sram_data_ok ? _GEN_9461 : _GEN_6389; // @[icache.scala 135:42]
  wire [184:0] _GEN_10486 = replace & io_inst_sram_data_ok ? _GEN_9462 : _GEN_6390; // @[icache.scala 135:42]
  wire [184:0] _GEN_10487 = replace & io_inst_sram_data_ok ? _GEN_9463 : _GEN_6391; // @[icache.scala 135:42]
  wire [184:0] _GEN_10488 = replace & io_inst_sram_data_ok ? _GEN_9464 : _GEN_6392; // @[icache.scala 135:42]
  wire [184:0] _GEN_10489 = replace & io_inst_sram_data_ok ? _GEN_9465 : _GEN_6393; // @[icache.scala 135:42]
  wire [184:0] _GEN_10490 = replace & io_inst_sram_data_ok ? _GEN_9466 : _GEN_6394; // @[icache.scala 135:42]
  wire [184:0] _GEN_10491 = replace & io_inst_sram_data_ok ? _GEN_9467 : _GEN_6395; // @[icache.scala 135:42]
  wire [184:0] _GEN_10492 = replace & io_inst_sram_data_ok ? _GEN_9468 : _GEN_6396; // @[icache.scala 135:42]
  wire [184:0] _GEN_10493 = replace & io_inst_sram_data_ok ? _GEN_9469 : _GEN_6397; // @[icache.scala 135:42]
  wire [184:0] _GEN_10494 = replace & io_inst_sram_data_ok ? _GEN_9470 : _GEN_6398; // @[icache.scala 135:42]
  wire [184:0] _GEN_10495 = replace & io_inst_sram_data_ok ? _GEN_9471 : _GEN_6399; // @[icache.scala 135:42]
  wire [184:0] _GEN_10496 = replace & io_inst_sram_data_ok ? _GEN_9472 : _GEN_6400; // @[icache.scala 135:42]
  wire [184:0] _GEN_10497 = replace & io_inst_sram_data_ok ? _GEN_9473 : _GEN_6401; // @[icache.scala 135:42]
  wire [184:0] _GEN_10498 = replace & io_inst_sram_data_ok ? _GEN_9474 : _GEN_6402; // @[icache.scala 135:42]
  wire [184:0] _GEN_10499 = replace & io_inst_sram_data_ok ? _GEN_9475 : _GEN_6403; // @[icache.scala 135:42]
  wire [184:0] _GEN_10500 = replace & io_inst_sram_data_ok ? _GEN_9476 : _GEN_6404; // @[icache.scala 135:42]
  wire [184:0] _GEN_10501 = replace & io_inst_sram_data_ok ? _GEN_9477 : _GEN_6405; // @[icache.scala 135:42]
  wire [184:0] _GEN_10502 = replace & io_inst_sram_data_ok ? _GEN_9478 : _GEN_6406; // @[icache.scala 135:42]
  wire [184:0] _GEN_10503 = replace & io_inst_sram_data_ok ? _GEN_9479 : _GEN_6407; // @[icache.scala 135:42]
  wire [184:0] _GEN_10504 = replace & io_inst_sram_data_ok ? _GEN_9480 : _GEN_6408; // @[icache.scala 135:42]
  wire [184:0] _GEN_10505 = replace & io_inst_sram_data_ok ? _GEN_9481 : _GEN_6409; // @[icache.scala 135:42]
  wire [184:0] _GEN_10506 = replace & io_inst_sram_data_ok ? _GEN_9482 : _GEN_6410; // @[icache.scala 135:42]
  wire [184:0] _GEN_10507 = replace & io_inst_sram_data_ok ? _GEN_9483 : _GEN_6411; // @[icache.scala 135:42]
  wire [184:0] _GEN_10508 = replace & io_inst_sram_data_ok ? _GEN_9484 : _GEN_6412; // @[icache.scala 135:42]
  wire [184:0] _GEN_10509 = replace & io_inst_sram_data_ok ? _GEN_9485 : _GEN_6413; // @[icache.scala 135:42]
  wire [184:0] _GEN_10510 = replace & io_inst_sram_data_ok ? _GEN_9486 : _GEN_6414; // @[icache.scala 135:42]
  wire [184:0] _GEN_10511 = replace & io_inst_sram_data_ok ? _GEN_9487 : _GEN_6415; // @[icache.scala 135:42]
  wire [184:0] _GEN_10512 = replace & io_inst_sram_data_ok ? _GEN_9488 : _GEN_6416; // @[icache.scala 135:42]
  wire [184:0] _GEN_10513 = replace & io_inst_sram_data_ok ? _GEN_9489 : _GEN_6417; // @[icache.scala 135:42]
  wire [184:0] _GEN_10514 = replace & io_inst_sram_data_ok ? _GEN_9490 : _GEN_6418; // @[icache.scala 135:42]
  wire [184:0] _GEN_10515 = replace & io_inst_sram_data_ok ? _GEN_9491 : _GEN_6419; // @[icache.scala 135:42]
  wire [184:0] _GEN_10516 = replace & io_inst_sram_data_ok ? _GEN_9492 : _GEN_6420; // @[icache.scala 135:42]
  wire [184:0] _GEN_10517 = replace & io_inst_sram_data_ok ? _GEN_9493 : _GEN_6421; // @[icache.scala 135:42]
  wire [184:0] _GEN_10518 = replace & io_inst_sram_data_ok ? _GEN_9494 : _GEN_6422; // @[icache.scala 135:42]
  wire [184:0] _GEN_10519 = replace & io_inst_sram_data_ok ? _GEN_9495 : _GEN_6423; // @[icache.scala 135:42]
  wire [184:0] _GEN_10520 = replace & io_inst_sram_data_ok ? _GEN_9496 : _GEN_6424; // @[icache.scala 135:42]
  wire [184:0] _GEN_10521 = replace & io_inst_sram_data_ok ? _GEN_9497 : _GEN_6425; // @[icache.scala 135:42]
  wire [184:0] _GEN_10522 = replace & io_inst_sram_data_ok ? _GEN_9498 : _GEN_6426; // @[icache.scala 135:42]
  wire [184:0] _GEN_10523 = replace & io_inst_sram_data_ok ? _GEN_9499 : _GEN_6427; // @[icache.scala 135:42]
  wire [184:0] _GEN_10524 = replace & io_inst_sram_data_ok ? _GEN_9500 : _GEN_6428; // @[icache.scala 135:42]
  wire [184:0] _GEN_10525 = replace & io_inst_sram_data_ok ? _GEN_9501 : _GEN_6429; // @[icache.scala 135:42]
  wire [184:0] _GEN_10526 = replace & io_inst_sram_data_ok ? _GEN_9502 : _GEN_6430; // @[icache.scala 135:42]
  wire [184:0] _GEN_10527 = replace & io_inst_sram_data_ok ? _GEN_9503 : _GEN_6431; // @[icache.scala 135:42]
  wire [184:0] _GEN_10528 = replace & io_inst_sram_data_ok ? _GEN_9504 : _GEN_6432; // @[icache.scala 135:42]
  wire [184:0] _GEN_10529 = replace & io_inst_sram_data_ok ? _GEN_9505 : _GEN_6433; // @[icache.scala 135:42]
  wire [184:0] _GEN_10530 = replace & io_inst_sram_data_ok ? _GEN_9506 : _GEN_6434; // @[icache.scala 135:42]
  wire [184:0] _GEN_10531 = replace & io_inst_sram_data_ok ? _GEN_9507 : _GEN_6435; // @[icache.scala 135:42]
  wire [184:0] _GEN_10532 = replace & io_inst_sram_data_ok ? _GEN_9508 : _GEN_6436; // @[icache.scala 135:42]
  wire [184:0] _GEN_10533 = replace & io_inst_sram_data_ok ? _GEN_9509 : _GEN_6437; // @[icache.scala 135:42]
  wire [184:0] _GEN_10534 = replace & io_inst_sram_data_ok ? _GEN_9510 : _GEN_6438; // @[icache.scala 135:42]
  wire [184:0] _GEN_10535 = replace & io_inst_sram_data_ok ? _GEN_9511 : _GEN_6439; // @[icache.scala 135:42]
  wire [184:0] _GEN_10536 = replace & io_inst_sram_data_ok ? _GEN_9512 : _GEN_6440; // @[icache.scala 135:42]
  wire [184:0] _GEN_10537 = replace & io_inst_sram_data_ok ? _GEN_9513 : _GEN_6441; // @[icache.scala 135:42]
  wire [184:0] _GEN_10538 = replace & io_inst_sram_data_ok ? _GEN_9514 : _GEN_6442; // @[icache.scala 135:42]
  wire [184:0] _GEN_10539 = replace & io_inst_sram_data_ok ? _GEN_9515 : _GEN_6443; // @[icache.scala 135:42]
  wire [184:0] _GEN_10540 = replace & io_inst_sram_data_ok ? _GEN_9516 : _GEN_6444; // @[icache.scala 135:42]
  wire [184:0] _GEN_10541 = replace & io_inst_sram_data_ok ? _GEN_9517 : _GEN_6445; // @[icache.scala 135:42]
  wire [184:0] _GEN_10542 = replace & io_inst_sram_data_ok ? _GEN_9518 : _GEN_6446; // @[icache.scala 135:42]
  wire [184:0] _GEN_10543 = replace & io_inst_sram_data_ok ? _GEN_9519 : _GEN_6447; // @[icache.scala 135:42]
  wire [184:0] _GEN_10544 = replace & io_inst_sram_data_ok ? _GEN_9520 : _GEN_6448; // @[icache.scala 135:42]
  wire [184:0] _GEN_10545 = replace & io_inst_sram_data_ok ? _GEN_9521 : _GEN_6449; // @[icache.scala 135:42]
  wire [184:0] _GEN_10546 = replace & io_inst_sram_data_ok ? _GEN_9522 : _GEN_6450; // @[icache.scala 135:42]
  wire [184:0] _GEN_10547 = replace & io_inst_sram_data_ok ? _GEN_9523 : _GEN_6451; // @[icache.scala 135:42]
  wire [184:0] _GEN_10548 = replace & io_inst_sram_data_ok ? _GEN_9524 : _GEN_6452; // @[icache.scala 135:42]
  wire [184:0] _GEN_10549 = replace & io_inst_sram_data_ok ? _GEN_9525 : _GEN_6453; // @[icache.scala 135:42]
  wire [184:0] _GEN_10550 = replace & io_inst_sram_data_ok ? _GEN_9526 : _GEN_6454; // @[icache.scala 135:42]
  wire [184:0] _GEN_10551 = replace & io_inst_sram_data_ok ? _GEN_9527 : _GEN_6455; // @[icache.scala 135:42]
  wire [184:0] _GEN_10552 = replace & io_inst_sram_data_ok ? _GEN_9528 : _GEN_6456; // @[icache.scala 135:42]
  wire [184:0] _GEN_10553 = replace & io_inst_sram_data_ok ? _GEN_9529 : _GEN_6457; // @[icache.scala 135:42]
  wire [184:0] _GEN_10554 = replace & io_inst_sram_data_ok ? _GEN_9530 : _GEN_6458; // @[icache.scala 135:42]
  wire [184:0] _GEN_10555 = replace & io_inst_sram_data_ok ? _GEN_9531 : _GEN_6459; // @[icache.scala 135:42]
  wire [184:0] _GEN_10556 = replace & io_inst_sram_data_ok ? _GEN_9532 : _GEN_6460; // @[icache.scala 135:42]
  wire [184:0] _GEN_10557 = replace & io_inst_sram_data_ok ? _GEN_9533 : _GEN_6461; // @[icache.scala 135:42]
  wire [184:0] _GEN_10558 = replace & io_inst_sram_data_ok ? _GEN_9534 : _GEN_6462; // @[icache.scala 135:42]
  wire [184:0] _GEN_10559 = replace & io_inst_sram_data_ok ? _GEN_9535 : _GEN_6463; // @[icache.scala 135:42]
  wire [184:0] _GEN_10560 = replace & io_inst_sram_data_ok ? _GEN_9536 : _GEN_6464; // @[icache.scala 135:42]
  wire [184:0] _GEN_10561 = replace & io_inst_sram_data_ok ? _GEN_9537 : _GEN_6465; // @[icache.scala 135:42]
  wire [184:0] _GEN_10562 = replace & io_inst_sram_data_ok ? _GEN_9538 : _GEN_6466; // @[icache.scala 135:42]
  wire [184:0] _GEN_10563 = replace & io_inst_sram_data_ok ? _GEN_9539 : _GEN_6467; // @[icache.scala 135:42]
  wire [184:0] _GEN_10564 = replace & io_inst_sram_data_ok ? _GEN_9540 : _GEN_6468; // @[icache.scala 135:42]
  wire [184:0] _GEN_10565 = replace & io_inst_sram_data_ok ? _GEN_9541 : _GEN_6469; // @[icache.scala 135:42]
  wire [184:0] _GEN_10566 = replace & io_inst_sram_data_ok ? _GEN_9542 : _GEN_6470; // @[icache.scala 135:42]
  wire [184:0] _GEN_10567 = replace & io_inst_sram_data_ok ? _GEN_9543 : _GEN_6471; // @[icache.scala 135:42]
  wire [184:0] _GEN_10568 = replace & io_inst_sram_data_ok ? _GEN_9544 : _GEN_6472; // @[icache.scala 135:42]
  wire [184:0] _GEN_10569 = replace & io_inst_sram_data_ok ? _GEN_9545 : _GEN_6473; // @[icache.scala 135:42]
  wire [184:0] _GEN_10570 = replace & io_inst_sram_data_ok ? _GEN_9546 : _GEN_6474; // @[icache.scala 135:42]
  wire [184:0] _GEN_10571 = replace & io_inst_sram_data_ok ? _GEN_9547 : _GEN_6475; // @[icache.scala 135:42]
  wire [184:0] _GEN_10572 = replace & io_inst_sram_data_ok ? _GEN_9548 : _GEN_6476; // @[icache.scala 135:42]
  wire [184:0] _GEN_10573 = replace & io_inst_sram_data_ok ? _GEN_9549 : _GEN_6477; // @[icache.scala 135:42]
  wire [184:0] _GEN_10574 = replace & io_inst_sram_data_ok ? _GEN_9550 : _GEN_6478; // @[icache.scala 135:42]
  wire [184:0] _GEN_10575 = replace & io_inst_sram_data_ok ? _GEN_9551 : _GEN_6479; // @[icache.scala 135:42]
  wire [184:0] _GEN_10576 = replace & io_inst_sram_data_ok ? _GEN_9552 : _GEN_6480; // @[icache.scala 135:42]
  wire [184:0] _GEN_10577 = replace & io_inst_sram_data_ok ? _GEN_9553 : _GEN_6481; // @[icache.scala 135:42]
  wire [184:0] _GEN_10578 = replace & io_inst_sram_data_ok ? _GEN_9554 : _GEN_6482; // @[icache.scala 135:42]
  wire [184:0] _GEN_10579 = replace & io_inst_sram_data_ok ? _GEN_9555 : _GEN_6483; // @[icache.scala 135:42]
  wire [184:0] _GEN_10580 = replace & io_inst_sram_data_ok ? _GEN_9556 : _GEN_6484; // @[icache.scala 135:42]
  wire [184:0] _GEN_10581 = replace & io_inst_sram_data_ok ? _GEN_9557 : _GEN_6485; // @[icache.scala 135:42]
  wire [184:0] _GEN_10582 = replace & io_inst_sram_data_ok ? _GEN_9558 : _GEN_6486; // @[icache.scala 135:42]
  wire [184:0] _GEN_10583 = replace & io_inst_sram_data_ok ? _GEN_9559 : _GEN_6487; // @[icache.scala 135:42]
  wire [184:0] _GEN_10584 = replace & io_inst_sram_data_ok ? _GEN_9560 : _GEN_6488; // @[icache.scala 135:42]
  wire [184:0] _GEN_10585 = replace & io_inst_sram_data_ok ? _GEN_9561 : _GEN_6489; // @[icache.scala 135:42]
  wire [184:0] _GEN_10586 = replace & io_inst_sram_data_ok ? _GEN_9562 : _GEN_6490; // @[icache.scala 135:42]
  wire [184:0] _GEN_10587 = replace & io_inst_sram_data_ok ? _GEN_9563 : _GEN_6491; // @[icache.scala 135:42]
  wire [184:0] _GEN_10588 = replace & io_inst_sram_data_ok ? _GEN_9564 : _GEN_6492; // @[icache.scala 135:42]
  wire [184:0] _GEN_10589 = replace & io_inst_sram_data_ok ? _GEN_9565 : _GEN_6493; // @[icache.scala 135:42]
  wire [184:0] _GEN_10590 = replace & io_inst_sram_data_ok ? _GEN_9566 : _GEN_6494; // @[icache.scala 135:42]
  wire [184:0] _GEN_10591 = replace & io_inst_sram_data_ok ? _GEN_9567 : _GEN_6495; // @[icache.scala 135:42]
  wire [184:0] _GEN_10592 = replace & io_inst_sram_data_ok ? _GEN_9568 : _GEN_6496; // @[icache.scala 135:42]
  wire [184:0] _GEN_10593 = replace & io_inst_sram_data_ok ? _GEN_9569 : _GEN_6497; // @[icache.scala 135:42]
  wire [184:0] _GEN_10594 = replace & io_inst_sram_data_ok ? _GEN_9570 : _GEN_6498; // @[icache.scala 135:42]
  wire [184:0] _GEN_10595 = replace & io_inst_sram_data_ok ? _GEN_9571 : _GEN_6499; // @[icache.scala 135:42]
  wire [184:0] _GEN_10596 = replace & io_inst_sram_data_ok ? _GEN_9572 : _GEN_6500; // @[icache.scala 135:42]
  wire [184:0] _GEN_10597 = replace & io_inst_sram_data_ok ? _GEN_9573 : _GEN_6501; // @[icache.scala 135:42]
  wire [184:0] _GEN_10598 = replace & io_inst_sram_data_ok ? _GEN_9574 : _GEN_6502; // @[icache.scala 135:42]
  wire [184:0] _GEN_10599 = replace & io_inst_sram_data_ok ? _GEN_9575 : _GEN_6503; // @[icache.scala 135:42]
  wire [184:0] _GEN_10600 = replace & io_inst_sram_data_ok ? _GEN_9576 : _GEN_6504; // @[icache.scala 135:42]
  wire [184:0] _GEN_10601 = replace & io_inst_sram_data_ok ? _GEN_9577 : _GEN_6505; // @[icache.scala 135:42]
  wire [184:0] _GEN_10602 = replace & io_inst_sram_data_ok ? _GEN_9578 : _GEN_6506; // @[icache.scala 135:42]
  wire [184:0] _GEN_10603 = replace & io_inst_sram_data_ok ? _GEN_9579 : _GEN_6507; // @[icache.scala 135:42]
  wire [184:0] _GEN_10604 = replace & io_inst_sram_data_ok ? _GEN_9580 : _GEN_6508; // @[icache.scala 135:42]
  wire [184:0] _GEN_10605 = replace & io_inst_sram_data_ok ? _GEN_9581 : _GEN_6509; // @[icache.scala 135:42]
  wire [184:0] _GEN_10606 = replace & io_inst_sram_data_ok ? _GEN_9582 : _GEN_6510; // @[icache.scala 135:42]
  wire [184:0] _GEN_10607 = replace & io_inst_sram_data_ok ? _GEN_9583 : _GEN_6511; // @[icache.scala 135:42]
  wire [184:0] _GEN_10608 = replace & io_inst_sram_data_ok ? _GEN_9584 : _GEN_6512; // @[icache.scala 135:42]
  wire [184:0] _GEN_10609 = replace & io_inst_sram_data_ok ? _GEN_9585 : _GEN_6513; // @[icache.scala 135:42]
  wire [184:0] _GEN_10610 = replace & io_inst_sram_data_ok ? _GEN_9586 : _GEN_6514; // @[icache.scala 135:42]
  wire [184:0] _GEN_10611 = replace & io_inst_sram_data_ok ? _GEN_9587 : _GEN_6515; // @[icache.scala 135:42]
  wire [184:0] _GEN_10612 = replace & io_inst_sram_data_ok ? _GEN_9588 : _GEN_6516; // @[icache.scala 135:42]
  wire [184:0] _GEN_10613 = replace & io_inst_sram_data_ok ? _GEN_9589 : _GEN_6517; // @[icache.scala 135:42]
  wire [184:0] _GEN_10614 = replace & io_inst_sram_data_ok ? _GEN_9590 : _GEN_6518; // @[icache.scala 135:42]
  wire [184:0] _GEN_10615 = replace & io_inst_sram_data_ok ? _GEN_9591 : _GEN_6519; // @[icache.scala 135:42]
  wire [184:0] _GEN_10616 = replace & io_inst_sram_data_ok ? _GEN_9592 : _GEN_6520; // @[icache.scala 135:42]
  wire [184:0] _GEN_10617 = replace & io_inst_sram_data_ok ? _GEN_9593 : _GEN_6521; // @[icache.scala 135:42]
  wire [184:0] _GEN_10618 = replace & io_inst_sram_data_ok ? _GEN_9594 : _GEN_6522; // @[icache.scala 135:42]
  wire [184:0] _GEN_10619 = replace & io_inst_sram_data_ok ? _GEN_9595 : _GEN_6523; // @[icache.scala 135:42]
  wire [184:0] _GEN_10620 = replace & io_inst_sram_data_ok ? _GEN_9596 : _GEN_6524; // @[icache.scala 135:42]
  wire [184:0] _GEN_10621 = replace & io_inst_sram_data_ok ? _GEN_9597 : _GEN_6525; // @[icache.scala 135:42]
  wire [184:0] _GEN_10622 = replace & io_inst_sram_data_ok ? _GEN_9598 : _GEN_6526; // @[icache.scala 135:42]
  wire [184:0] _GEN_10623 = replace & io_inst_sram_data_ok ? _GEN_9599 : _GEN_6527; // @[icache.scala 135:42]
  wire [184:0] _GEN_10624 = replace & io_inst_sram_data_ok ? _GEN_9600 : _GEN_6528; // @[icache.scala 135:42]
  wire [184:0] _GEN_10625 = replace & io_inst_sram_data_ok ? _GEN_9601 : _GEN_6529; // @[icache.scala 135:42]
  wire [184:0] _GEN_10626 = replace & io_inst_sram_data_ok ? _GEN_9602 : _GEN_6530; // @[icache.scala 135:42]
  wire [184:0] _GEN_10627 = replace & io_inst_sram_data_ok ? _GEN_9603 : _GEN_6531; // @[icache.scala 135:42]
  wire [184:0] _GEN_10628 = replace & io_inst_sram_data_ok ? _GEN_9604 : _GEN_6532; // @[icache.scala 135:42]
  wire [184:0] _GEN_10629 = replace & io_inst_sram_data_ok ? _GEN_9605 : _GEN_6533; // @[icache.scala 135:42]
  wire [184:0] _GEN_10630 = replace & io_inst_sram_data_ok ? _GEN_9606 : _GEN_6534; // @[icache.scala 135:42]
  wire [184:0] _GEN_10631 = replace & io_inst_sram_data_ok ? _GEN_9607 : _GEN_6535; // @[icache.scala 135:42]
  wire [184:0] _GEN_10632 = replace & io_inst_sram_data_ok ? _GEN_9608 : _GEN_6536; // @[icache.scala 135:42]
  wire [184:0] _GEN_10633 = replace & io_inst_sram_data_ok ? _GEN_9609 : _GEN_6537; // @[icache.scala 135:42]
  wire [184:0] _GEN_10634 = replace & io_inst_sram_data_ok ? _GEN_9610 : _GEN_6538; // @[icache.scala 135:42]
  wire [184:0] _GEN_10635 = replace & io_inst_sram_data_ok ? _GEN_9611 : _GEN_6539; // @[icache.scala 135:42]
  wire [184:0] _GEN_10636 = replace & io_inst_sram_data_ok ? _GEN_9612 : _GEN_6540; // @[icache.scala 135:42]
  wire [184:0] _GEN_10637 = replace & io_inst_sram_data_ok ? _GEN_9613 : _GEN_6541; // @[icache.scala 135:42]
  wire [184:0] _GEN_10638 = replace & io_inst_sram_data_ok ? _GEN_9614 : _GEN_6542; // @[icache.scala 135:42]
  wire [184:0] _GEN_10639 = replace & io_inst_sram_data_ok ? _GEN_9615 : _GEN_6543; // @[icache.scala 135:42]
  wire [184:0] _GEN_10640 = replace & io_inst_sram_data_ok ? _GEN_9616 : _GEN_6544; // @[icache.scala 135:42]
  wire [184:0] _GEN_10641 = replace & io_inst_sram_data_ok ? _GEN_9617 : _GEN_6545; // @[icache.scala 135:42]
  wire [184:0] _GEN_10642 = replace & io_inst_sram_data_ok ? _GEN_9618 : _GEN_6546; // @[icache.scala 135:42]
  wire [184:0] _GEN_10643 = replace & io_inst_sram_data_ok ? _GEN_9619 : _GEN_6547; // @[icache.scala 135:42]
  wire [184:0] _GEN_10644 = replace & io_inst_sram_data_ok ? _GEN_9620 : _GEN_6548; // @[icache.scala 135:42]
  wire [184:0] _GEN_10645 = replace & io_inst_sram_data_ok ? _GEN_9621 : _GEN_6549; // @[icache.scala 135:42]
  wire [184:0] _GEN_10646 = replace & io_inst_sram_data_ok ? _GEN_9622 : _GEN_6550; // @[icache.scala 135:42]
  wire [184:0] _GEN_10647 = replace & io_inst_sram_data_ok ? _GEN_9623 : _GEN_6551; // @[icache.scala 135:42]
  wire [184:0] _GEN_10648 = replace & io_inst_sram_data_ok ? _GEN_9624 : _GEN_6552; // @[icache.scala 135:42]
  wire [184:0] _GEN_10649 = replace & io_inst_sram_data_ok ? _GEN_9625 : _GEN_6553; // @[icache.scala 135:42]
  wire [184:0] _GEN_10650 = replace & io_inst_sram_data_ok ? _GEN_9626 : _GEN_6554; // @[icache.scala 135:42]
  wire [184:0] _GEN_10651 = replace & io_inst_sram_data_ok ? _GEN_9627 : _GEN_6555; // @[icache.scala 135:42]
  wire [184:0] _GEN_10652 = replace & io_inst_sram_data_ok ? _GEN_9628 : _GEN_6556; // @[icache.scala 135:42]
  wire [184:0] _GEN_10653 = replace & io_inst_sram_data_ok ? _GEN_9629 : _GEN_6557; // @[icache.scala 135:42]
  wire [184:0] _GEN_10654 = replace & io_inst_sram_data_ok ? _GEN_9630 : _GEN_6558; // @[icache.scala 135:42]
  wire [184:0] _GEN_10655 = replace & io_inst_sram_data_ok ? _GEN_9631 : _GEN_6559; // @[icache.scala 135:42]
  wire [184:0] _GEN_10656 = replace & io_inst_sram_data_ok ? _GEN_9632 : _GEN_6560; // @[icache.scala 135:42]
  wire [184:0] _GEN_10657 = replace & io_inst_sram_data_ok ? _GEN_9633 : _GEN_6561; // @[icache.scala 135:42]
  wire [184:0] _GEN_10658 = replace & io_inst_sram_data_ok ? _GEN_9634 : _GEN_6562; // @[icache.scala 135:42]
  wire [184:0] _GEN_10659 = replace & io_inst_sram_data_ok ? _GEN_9635 : _GEN_6563; // @[icache.scala 135:42]
  wire [184:0] _GEN_10660 = replace & io_inst_sram_data_ok ? _GEN_9636 : _GEN_6564; // @[icache.scala 135:42]
  wire [184:0] _GEN_10661 = replace & io_inst_sram_data_ok ? _GEN_9637 : _GEN_6565; // @[icache.scala 135:42]
  wire [184:0] _GEN_10662 = replace & io_inst_sram_data_ok ? _GEN_9638 : _GEN_6566; // @[icache.scala 135:42]
  wire [184:0] _GEN_10663 = replace & io_inst_sram_data_ok ? _GEN_9639 : _GEN_6567; // @[icache.scala 135:42]
  wire [184:0] _GEN_10664 = replace & io_inst_sram_data_ok ? _GEN_9640 : _GEN_6568; // @[icache.scala 135:42]
  wire [184:0] _GEN_10665 = replace & io_inst_sram_data_ok ? _GEN_9641 : _GEN_6569; // @[icache.scala 135:42]
  wire [184:0] _GEN_10666 = replace & io_inst_sram_data_ok ? _GEN_9642 : _GEN_6570; // @[icache.scala 135:42]
  wire [184:0] _GEN_10667 = replace & io_inst_sram_data_ok ? _GEN_9643 : _GEN_6571; // @[icache.scala 135:42]
  wire [184:0] _GEN_10668 = replace & io_inst_sram_data_ok ? _GEN_9644 : _GEN_6572; // @[icache.scala 135:42]
  wire [184:0] _GEN_10669 = replace & io_inst_sram_data_ok ? _GEN_9645 : _GEN_6573; // @[icache.scala 135:42]
  wire [184:0] _GEN_10670 = replace & io_inst_sram_data_ok ? _GEN_9646 : _GEN_6574; // @[icache.scala 135:42]
  wire [184:0] _GEN_10671 = replace & io_inst_sram_data_ok ? _GEN_9647 : _GEN_6575; // @[icache.scala 135:42]
  wire [184:0] _GEN_10672 = replace & io_inst_sram_data_ok ? _GEN_9648 : _GEN_6576; // @[icache.scala 135:42]
  wire [184:0] _GEN_10673 = replace & io_inst_sram_data_ok ? _GEN_9649 : _GEN_6577; // @[icache.scala 135:42]
  wire [184:0] _GEN_10674 = replace & io_inst_sram_data_ok ? _GEN_9650 : _GEN_6578; // @[icache.scala 135:42]
  wire [184:0] _GEN_10675 = replace & io_inst_sram_data_ok ? _GEN_9651 : _GEN_6579; // @[icache.scala 135:42]
  wire [184:0] _GEN_10676 = replace & io_inst_sram_data_ok ? _GEN_9652 : _GEN_6580; // @[icache.scala 135:42]
  wire [184:0] _GEN_10677 = replace & io_inst_sram_data_ok ? _GEN_9653 : _GEN_6581; // @[icache.scala 135:42]
  wire [184:0] _GEN_10678 = replace & io_inst_sram_data_ok ? _GEN_9654 : _GEN_6582; // @[icache.scala 135:42]
  wire [184:0] _GEN_10679 = replace & io_inst_sram_data_ok ? _GEN_9655 : _GEN_6583; // @[icache.scala 135:42]
  wire [184:0] _GEN_10680 = replace & io_inst_sram_data_ok ? _GEN_9656 : _GEN_6584; // @[icache.scala 135:42]
  wire [184:0] _GEN_10681 = replace & io_inst_sram_data_ok ? _GEN_9657 : _GEN_6585; // @[icache.scala 135:42]
  wire [184:0] _GEN_10682 = replace & io_inst_sram_data_ok ? _GEN_9658 : _GEN_6586; // @[icache.scala 135:42]
  wire [184:0] _GEN_10683 = replace & io_inst_sram_data_ok ? _GEN_9659 : _GEN_6587; // @[icache.scala 135:42]
  wire [184:0] _GEN_10684 = replace & io_inst_sram_data_ok ? _GEN_9660 : _GEN_6588; // @[icache.scala 135:42]
  wire [184:0] _GEN_10685 = replace & io_inst_sram_data_ok ? _GEN_9661 : _GEN_6589; // @[icache.scala 135:42]
  wire [184:0] _GEN_10686 = replace & io_inst_sram_data_ok ? _GEN_9662 : _GEN_6590; // @[icache.scala 135:42]
  wire [184:0] _GEN_10687 = replace & io_inst_sram_data_ok ? _GEN_9663 : _GEN_6591; // @[icache.scala 135:42]
  wire [184:0] _GEN_10688 = replace & io_inst_sram_data_ok ? _GEN_9664 : _GEN_6592; // @[icache.scala 135:42]
  wire [184:0] _GEN_10689 = replace & io_inst_sram_data_ok ? _GEN_9665 : _GEN_6593; // @[icache.scala 135:42]
  wire [184:0] _GEN_10690 = replace & io_inst_sram_data_ok ? _GEN_9666 : _GEN_6594; // @[icache.scala 135:42]
  wire [184:0] _GEN_10691 = replace & io_inst_sram_data_ok ? _GEN_9667 : _GEN_6595; // @[icache.scala 135:42]
  wire [184:0] _GEN_10692 = replace & io_inst_sram_data_ok ? _GEN_9668 : _GEN_6596; // @[icache.scala 135:42]
  wire [184:0] _GEN_10693 = replace & io_inst_sram_data_ok ? _GEN_9669 : _GEN_6597; // @[icache.scala 135:42]
  wire [184:0] _GEN_10694 = replace & io_inst_sram_data_ok ? _GEN_9670 : _GEN_6598; // @[icache.scala 135:42]
  wire [184:0] _GEN_10695 = replace & io_inst_sram_data_ok ? _GEN_9671 : _GEN_6599; // @[icache.scala 135:42]
  wire [184:0] _GEN_10696 = replace & io_inst_sram_data_ok ? _GEN_9672 : _GEN_6600; // @[icache.scala 135:42]
  wire [184:0] _GEN_10697 = replace & io_inst_sram_data_ok ? _GEN_9673 : _GEN_6601; // @[icache.scala 135:42]
  wire [184:0] _GEN_10698 = replace & io_inst_sram_data_ok ? _GEN_9674 : _GEN_6602; // @[icache.scala 135:42]
  wire [184:0] _GEN_10699 = replace & io_inst_sram_data_ok ? _GEN_9675 : _GEN_6603; // @[icache.scala 135:42]
  wire [184:0] _GEN_10700 = replace & io_inst_sram_data_ok ? _GEN_9676 : _GEN_6604; // @[icache.scala 135:42]
  wire [184:0] _GEN_10701 = replace & io_inst_sram_data_ok ? _GEN_9677 : _GEN_6605; // @[icache.scala 135:42]
  wire [184:0] _GEN_10702 = replace & io_inst_sram_data_ok ? _GEN_9678 : _GEN_6606; // @[icache.scala 135:42]
  wire [184:0] _GEN_10703 = replace & io_inst_sram_data_ok ? _GEN_9679 : _GEN_6607; // @[icache.scala 135:42]
  wire [184:0] _GEN_10704 = replace & io_inst_sram_data_ok ? _GEN_9680 : _GEN_6608; // @[icache.scala 135:42]
  wire [184:0] _GEN_10705 = replace & io_inst_sram_data_ok ? _GEN_9681 : _GEN_6609; // @[icache.scala 135:42]
  wire [184:0] _GEN_10706 = replace & io_inst_sram_data_ok ? _GEN_9682 : _GEN_6610; // @[icache.scala 135:42]
  wire [184:0] _GEN_10707 = replace & io_inst_sram_data_ok ? _GEN_9683 : _GEN_6611; // @[icache.scala 135:42]
  wire [184:0] _GEN_10708 = replace & io_inst_sram_data_ok ? _GEN_9684 : _GEN_6612; // @[icache.scala 135:42]
  wire [184:0] _GEN_10709 = replace & io_inst_sram_data_ok ? _GEN_9685 : _GEN_6613; // @[icache.scala 135:42]
  wire [184:0] _GEN_10710 = replace & io_inst_sram_data_ok ? _GEN_9686 : _GEN_6614; // @[icache.scala 135:42]
  wire [184:0] _GEN_10711 = replace & io_inst_sram_data_ok ? _GEN_9687 : _GEN_6615; // @[icache.scala 135:42]
  wire [184:0] _GEN_10712 = replace & io_inst_sram_data_ok ? _GEN_9688 : _GEN_6616; // @[icache.scala 135:42]
  wire [184:0] _GEN_10713 = replace & io_inst_sram_data_ok ? _GEN_9689 : _GEN_6617; // @[icache.scala 135:42]
  wire [184:0] _GEN_10714 = replace & io_inst_sram_data_ok ? _GEN_9690 : _GEN_6618; // @[icache.scala 135:42]
  wire [184:0] _GEN_10715 = replace & io_inst_sram_data_ok ? _GEN_9691 : _GEN_6619; // @[icache.scala 135:42]
  wire [184:0] _GEN_10716 = replace & io_inst_sram_data_ok ? _GEN_9692 : _GEN_6620; // @[icache.scala 135:42]
  wire [184:0] _GEN_10717 = replace & io_inst_sram_data_ok ? _GEN_9693 : _GEN_6621; // @[icache.scala 135:42]
  wire [184:0] _GEN_10718 = replace & io_inst_sram_data_ok ? _GEN_9694 : _GEN_6622; // @[icache.scala 135:42]
  wire [184:0] _GEN_10719 = replace & io_inst_sram_data_ok ? _GEN_9695 : _GEN_6623; // @[icache.scala 135:42]
  wire [184:0] _GEN_10720 = replace & io_inst_sram_data_ok ? _GEN_9696 : _GEN_6624; // @[icache.scala 135:42]
  wire [184:0] _GEN_10721 = replace & io_inst_sram_data_ok ? _GEN_9697 : _GEN_6625; // @[icache.scala 135:42]
  wire [184:0] _GEN_10722 = replace & io_inst_sram_data_ok ? _GEN_9698 : _GEN_6626; // @[icache.scala 135:42]
  wire [184:0] _GEN_10723 = replace & io_inst_sram_data_ok ? _GEN_9699 : _GEN_6627; // @[icache.scala 135:42]
  wire [184:0] _GEN_10724 = replace & io_inst_sram_data_ok ? _GEN_9700 : _GEN_6628; // @[icache.scala 135:42]
  wire [184:0] _GEN_10725 = replace & io_inst_sram_data_ok ? _GEN_9701 : _GEN_6629; // @[icache.scala 135:42]
  wire [184:0] _GEN_10726 = replace & io_inst_sram_data_ok ? _GEN_9702 : _GEN_6630; // @[icache.scala 135:42]
  wire [184:0] _GEN_10727 = replace & io_inst_sram_data_ok ? _GEN_9703 : _GEN_6631; // @[icache.scala 135:42]
  wire [184:0] _GEN_10728 = replace & io_inst_sram_data_ok ? _GEN_9704 : _GEN_6632; // @[icache.scala 135:42]
  wire [184:0] _GEN_10729 = replace & io_inst_sram_data_ok ? _GEN_9705 : _GEN_6633; // @[icache.scala 135:42]
  wire [184:0] _GEN_10730 = replace & io_inst_sram_data_ok ? _GEN_9706 : _GEN_6634; // @[icache.scala 135:42]
  wire [184:0] _GEN_10731 = replace & io_inst_sram_data_ok ? _GEN_9707 : _GEN_6635; // @[icache.scala 135:42]
  wire [184:0] _GEN_10732 = replace & io_inst_sram_data_ok ? _GEN_9708 : _GEN_6636; // @[icache.scala 135:42]
  wire [184:0] _GEN_10733 = replace & io_inst_sram_data_ok ? _GEN_9709 : _GEN_6637; // @[icache.scala 135:42]
  wire [184:0] _GEN_10734 = replace & io_inst_sram_data_ok ? _GEN_9710 : _GEN_6638; // @[icache.scala 135:42]
  wire [184:0] _GEN_10735 = replace & io_inst_sram_data_ok ? _GEN_9711 : _GEN_6639; // @[icache.scala 135:42]
  wire [184:0] _GEN_10736 = replace & io_inst_sram_data_ok ? _GEN_9712 : _GEN_6640; // @[icache.scala 135:42]
  wire [184:0] _GEN_10737 = replace & io_inst_sram_data_ok ? _GEN_9713 : _GEN_6641; // @[icache.scala 135:42]
  wire [184:0] _GEN_10738 = replace & io_inst_sram_data_ok ? _GEN_9714 : _GEN_6642; // @[icache.scala 135:42]
  wire [184:0] _GEN_10739 = replace & io_inst_sram_data_ok ? _GEN_9715 : _GEN_6643; // @[icache.scala 135:42]
  wire [184:0] _GEN_10740 = replace & io_inst_sram_data_ok ? _GEN_9716 : _GEN_6644; // @[icache.scala 135:42]
  wire [184:0] _GEN_10741 = replace & io_inst_sram_data_ok ? _GEN_9717 : _GEN_6645; // @[icache.scala 135:42]
  wire [184:0] _GEN_10742 = replace & io_inst_sram_data_ok ? _GEN_9718 : _GEN_6646; // @[icache.scala 135:42]
  wire [184:0] _GEN_10743 = replace & io_inst_sram_data_ok ? _GEN_9719 : _GEN_6647; // @[icache.scala 135:42]
  wire [184:0] _GEN_10744 = replace & io_inst_sram_data_ok ? _GEN_9720 : _GEN_6648; // @[icache.scala 135:42]
  wire [184:0] _GEN_10745 = replace & io_inst_sram_data_ok ? _GEN_9721 : _GEN_6649; // @[icache.scala 135:42]
  wire [184:0] _GEN_10746 = replace & io_inst_sram_data_ok ? _GEN_9722 : _GEN_6650; // @[icache.scala 135:42]
  wire [184:0] _GEN_10747 = replace & io_inst_sram_data_ok ? _GEN_9723 : _GEN_6651; // @[icache.scala 135:42]
  wire [184:0] _GEN_10748 = replace & io_inst_sram_data_ok ? _GEN_9724 : _GEN_6652; // @[icache.scala 135:42]
  wire [184:0] _GEN_10749 = replace & io_inst_sram_data_ok ? _GEN_9725 : _GEN_6653; // @[icache.scala 135:42]
  wire [184:0] _GEN_10750 = replace & io_inst_sram_data_ok ? _GEN_9726 : _GEN_6654; // @[icache.scala 135:42]
  wire [184:0] _GEN_10751 = replace & io_inst_sram_data_ok ? _GEN_9727 : _GEN_6655; // @[icache.scala 135:42]
  wire [184:0] _GEN_10752 = replace & io_inst_sram_data_ok ? _GEN_9728 : _GEN_6656; // @[icache.scala 135:42]
  wire [184:0] _GEN_10753 = replace & io_inst_sram_data_ok ? _GEN_9729 : _GEN_6657; // @[icache.scala 135:42]
  wire [184:0] _GEN_10754 = replace & io_inst_sram_data_ok ? _GEN_9730 : _GEN_6658; // @[icache.scala 135:42]
  wire [184:0] _GEN_10755 = replace & io_inst_sram_data_ok ? _GEN_9731 : _GEN_6659; // @[icache.scala 135:42]
  wire [184:0] _GEN_10756 = replace & io_inst_sram_data_ok ? _GEN_9732 : _GEN_6660; // @[icache.scala 135:42]
  wire [184:0] _GEN_10757 = replace & io_inst_sram_data_ok ? _GEN_9733 : _GEN_6661; // @[icache.scala 135:42]
  wire [184:0] _GEN_10758 = replace & io_inst_sram_data_ok ? _GEN_9734 : _GEN_6662; // @[icache.scala 135:42]
  wire [184:0] _GEN_10759 = replace & io_inst_sram_data_ok ? _GEN_9735 : _GEN_6663; // @[icache.scala 135:42]
  wire [184:0] _GEN_10760 = replace & io_inst_sram_data_ok ? _GEN_9736 : _GEN_6664; // @[icache.scala 135:42]
  wire [184:0] _GEN_10761 = replace & io_inst_sram_data_ok ? _GEN_9737 : _GEN_6665; // @[icache.scala 135:42]
  wire [184:0] _GEN_10762 = replace & io_inst_sram_data_ok ? _GEN_9738 : _GEN_6666; // @[icache.scala 135:42]
  wire [184:0] _GEN_10763 = replace & io_inst_sram_data_ok ? _GEN_9739 : _GEN_6667; // @[icache.scala 135:42]
  wire [184:0] _GEN_10764 = replace & io_inst_sram_data_ok ? _GEN_9740 : _GEN_6668; // @[icache.scala 135:42]
  wire [184:0] _GEN_10765 = replace & io_inst_sram_data_ok ? _GEN_9741 : _GEN_6669; // @[icache.scala 135:42]
  wire [184:0] _GEN_10766 = replace & io_inst_sram_data_ok ? _GEN_9742 : _GEN_6670; // @[icache.scala 135:42]
  wire [184:0] _GEN_10767 = replace & io_inst_sram_data_ok ? _GEN_9743 : _GEN_6671; // @[icache.scala 135:42]
  wire [184:0] _GEN_10768 = replace & io_inst_sram_data_ok ? _GEN_9744 : _GEN_6672; // @[icache.scala 135:42]
  wire [184:0] _GEN_10769 = replace & io_inst_sram_data_ok ? _GEN_9745 : _GEN_6673; // @[icache.scala 135:42]
  wire [184:0] _GEN_10770 = replace & io_inst_sram_data_ok ? _GEN_9746 : _GEN_6674; // @[icache.scala 135:42]
  wire [184:0] _GEN_10771 = replace & io_inst_sram_data_ok ? _GEN_9747 : _GEN_6675; // @[icache.scala 135:42]
  wire [184:0] _GEN_10772 = replace & io_inst_sram_data_ok ? _GEN_9748 : _GEN_6676; // @[icache.scala 135:42]
  wire [184:0] _GEN_10773 = replace & io_inst_sram_data_ok ? _GEN_9749 : _GEN_6677; // @[icache.scala 135:42]
  wire [184:0] _GEN_10774 = replace & io_inst_sram_data_ok ? _GEN_9750 : _GEN_6678; // @[icache.scala 135:42]
  wire [184:0] _GEN_10775 = replace & io_inst_sram_data_ok ? _GEN_9751 : _GEN_6679; // @[icache.scala 135:42]
  wire [184:0] _GEN_10776 = replace & io_inst_sram_data_ok ? _GEN_9752 : _GEN_6680; // @[icache.scala 135:42]
  wire [184:0] _GEN_10777 = replace & io_inst_sram_data_ok ? _GEN_9753 : _GEN_6681; // @[icache.scala 135:42]
  wire [184:0] _GEN_10778 = replace & io_inst_sram_data_ok ? _GEN_9754 : _GEN_6682; // @[icache.scala 135:42]
  wire [184:0] _GEN_10779 = replace & io_inst_sram_data_ok ? _GEN_9755 : _GEN_6683; // @[icache.scala 135:42]
  wire [184:0] _GEN_10780 = replace & io_inst_sram_data_ok ? _GEN_9756 : _GEN_6684; // @[icache.scala 135:42]
  wire [184:0] _GEN_10781 = replace & io_inst_sram_data_ok ? _GEN_9757 : _GEN_6685; // @[icache.scala 135:42]
  wire [184:0] _GEN_10782 = replace & io_inst_sram_data_ok ? _GEN_9758 : _GEN_6686; // @[icache.scala 135:42]
  wire [184:0] _GEN_10783 = replace & io_inst_sram_data_ok ? _GEN_9759 : _GEN_6687; // @[icache.scala 135:42]
  wire [184:0] _GEN_10784 = replace & io_inst_sram_data_ok ? _GEN_9760 : _GEN_6688; // @[icache.scala 135:42]
  wire [184:0] _GEN_10785 = replace & io_inst_sram_data_ok ? _GEN_9761 : _GEN_6689; // @[icache.scala 135:42]
  wire [184:0] _GEN_10786 = replace & io_inst_sram_data_ok ? _GEN_9762 : _GEN_6690; // @[icache.scala 135:42]
  wire [184:0] _GEN_10787 = replace & io_inst_sram_data_ok ? _GEN_9763 : _GEN_6691; // @[icache.scala 135:42]
  wire [184:0] _GEN_10788 = replace & io_inst_sram_data_ok ? _GEN_9764 : _GEN_6692; // @[icache.scala 135:42]
  wire [184:0] _GEN_10789 = replace & io_inst_sram_data_ok ? _GEN_9765 : _GEN_6693; // @[icache.scala 135:42]
  wire [184:0] _GEN_10790 = replace & io_inst_sram_data_ok ? _GEN_9766 : _GEN_6694; // @[icache.scala 135:42]
  wire [184:0] _GEN_10791 = replace & io_inst_sram_data_ok ? _GEN_9767 : _GEN_6695; // @[icache.scala 135:42]
  wire [184:0] _GEN_10792 = replace & io_inst_sram_data_ok ? _GEN_9768 : _GEN_6696; // @[icache.scala 135:42]
  wire [184:0] _GEN_10793 = replace & io_inst_sram_data_ok ? _GEN_9769 : _GEN_6697; // @[icache.scala 135:42]
  wire [184:0] _GEN_10794 = replace & io_inst_sram_data_ok ? _GEN_9770 : _GEN_6698; // @[icache.scala 135:42]
  wire [184:0] _GEN_10795 = replace & io_inst_sram_data_ok ? _GEN_9771 : _GEN_6699; // @[icache.scala 135:42]
  wire [184:0] _GEN_10796 = replace & io_inst_sram_data_ok ? _GEN_9772 : _GEN_6700; // @[icache.scala 135:42]
  wire [184:0] _GEN_10797 = replace & io_inst_sram_data_ok ? _GEN_9773 : _GEN_6701; // @[icache.scala 135:42]
  wire [184:0] _GEN_10798 = replace & io_inst_sram_data_ok ? _GEN_9774 : _GEN_6702; // @[icache.scala 135:42]
  wire [184:0] _GEN_10799 = replace & io_inst_sram_data_ok ? _GEN_9775 : _GEN_6703; // @[icache.scala 135:42]
  wire [184:0] _GEN_10800 = replace & io_inst_sram_data_ok ? _GEN_9776 : _GEN_6704; // @[icache.scala 135:42]
  wire [184:0] _GEN_10801 = replace & io_inst_sram_data_ok ? _GEN_9777 : _GEN_6705; // @[icache.scala 135:42]
  wire [184:0] _GEN_10802 = replace & io_inst_sram_data_ok ? _GEN_9778 : _GEN_6706; // @[icache.scala 135:42]
  wire [184:0] _GEN_10803 = replace & io_inst_sram_data_ok ? _GEN_9779 : _GEN_6707; // @[icache.scala 135:42]
  wire [184:0] _GEN_10804 = replace & io_inst_sram_data_ok ? _GEN_9780 : _GEN_6708; // @[icache.scala 135:42]
  wire [184:0] _GEN_10805 = replace & io_inst_sram_data_ok ? _GEN_9781 : _GEN_6709; // @[icache.scala 135:42]
  wire [184:0] _GEN_10806 = replace & io_inst_sram_data_ok ? _GEN_9782 : _GEN_6710; // @[icache.scala 135:42]
  wire [184:0] _GEN_10807 = replace & io_inst_sram_data_ok ? _GEN_9783 : _GEN_6711; // @[icache.scala 135:42]
  wire [184:0] _GEN_10808 = replace & io_inst_sram_data_ok ? _GEN_9784 : _GEN_6712; // @[icache.scala 135:42]
  wire [184:0] _GEN_10809 = replace & io_inst_sram_data_ok ? _GEN_9785 : _GEN_6713; // @[icache.scala 135:42]
  wire [184:0] _GEN_10810 = replace & io_inst_sram_data_ok ? _GEN_9786 : _GEN_6714; // @[icache.scala 135:42]
  wire [184:0] _GEN_10811 = replace & io_inst_sram_data_ok ? _GEN_9787 : _GEN_6715; // @[icache.scala 135:42]
  wire [184:0] _GEN_10812 = replace & io_inst_sram_data_ok ? _GEN_9788 : _GEN_6716; // @[icache.scala 135:42]
  wire [184:0] _GEN_10813 = replace & io_inst_sram_data_ok ? _GEN_9789 : _GEN_6717; // @[icache.scala 135:42]
  wire [184:0] _GEN_10814 = replace & io_inst_sram_data_ok ? _GEN_9790 : _GEN_6718; // @[icache.scala 135:42]
  wire [184:0] _GEN_10815 = replace & io_inst_sram_data_ok ? _GEN_9791 : _GEN_6719; // @[icache.scala 135:42]
  wire [184:0] _GEN_10816 = replace & io_inst_sram_data_ok ? _GEN_9792 : _GEN_6720; // @[icache.scala 135:42]
  wire [184:0] _GEN_10817 = replace & io_inst_sram_data_ok ? _GEN_9793 : _GEN_6721; // @[icache.scala 135:42]
  wire [184:0] _GEN_10818 = replace & io_inst_sram_data_ok ? _GEN_9794 : _GEN_6722; // @[icache.scala 135:42]
  wire [184:0] _GEN_10819 = replace & io_inst_sram_data_ok ? _GEN_9795 : _GEN_6723; // @[icache.scala 135:42]
  wire [184:0] _GEN_10820 = replace & io_inst_sram_data_ok ? _GEN_9796 : _GEN_6724; // @[icache.scala 135:42]
  wire [184:0] _GEN_10821 = replace & io_inst_sram_data_ok ? _GEN_9797 : _GEN_6725; // @[icache.scala 135:42]
  wire [184:0] _GEN_10822 = replace & io_inst_sram_data_ok ? _GEN_9798 : _GEN_6726; // @[icache.scala 135:42]
  wire [184:0] _GEN_10823 = replace & io_inst_sram_data_ok ? _GEN_9799 : _GEN_6727; // @[icache.scala 135:42]
  wire [184:0] _GEN_10824 = replace & io_inst_sram_data_ok ? _GEN_9800 : _GEN_6728; // @[icache.scala 135:42]
  wire [184:0] _GEN_10825 = replace & io_inst_sram_data_ok ? _GEN_9801 : _GEN_6729; // @[icache.scala 135:42]
  wire [184:0] _GEN_10826 = replace & io_inst_sram_data_ok ? _GEN_9802 : _GEN_6730; // @[icache.scala 135:42]
  wire [184:0] _GEN_10827 = replace & io_inst_sram_data_ok ? _GEN_9803 : _GEN_6731; // @[icache.scala 135:42]
  wire [184:0] _GEN_10828 = replace & io_inst_sram_data_ok ? _GEN_9804 : _GEN_6732; // @[icache.scala 135:42]
  wire [184:0] _GEN_10829 = replace & io_inst_sram_data_ok ? _GEN_9805 : _GEN_6733; // @[icache.scala 135:42]
  wire [184:0] _GEN_10830 = replace & io_inst_sram_data_ok ? _GEN_9806 : _GEN_6734; // @[icache.scala 135:42]
  wire [184:0] _GEN_10831 = replace & io_inst_sram_data_ok ? _GEN_9807 : _GEN_6735; // @[icache.scala 135:42]
  wire [184:0] _GEN_10832 = replace & io_inst_sram_data_ok ? _GEN_9808 : _GEN_6736; // @[icache.scala 135:42]
  wire [184:0] _GEN_10833 = replace & io_inst_sram_data_ok ? _GEN_9809 : _GEN_6737; // @[icache.scala 135:42]
  wire [184:0] _GEN_10834 = replace & io_inst_sram_data_ok ? _GEN_9810 : _GEN_6738; // @[icache.scala 135:42]
  wire [184:0] _GEN_10835 = replace & io_inst_sram_data_ok ? _GEN_9811 : _GEN_6739; // @[icache.scala 135:42]
  wire [184:0] _GEN_10836 = replace & io_inst_sram_data_ok ? _GEN_9812 : _GEN_6740; // @[icache.scala 135:42]
  wire [184:0] _GEN_10837 = replace & io_inst_sram_data_ok ? _GEN_9813 : _GEN_6741; // @[icache.scala 135:42]
  wire [184:0] _GEN_10838 = replace & io_inst_sram_data_ok ? _GEN_9814 : _GEN_6742; // @[icache.scala 135:42]
  wire [184:0] _GEN_10839 = replace & io_inst_sram_data_ok ? _GEN_9815 : _GEN_6743; // @[icache.scala 135:42]
  wire [184:0] _GEN_10840 = replace & io_inst_sram_data_ok ? _GEN_9816 : _GEN_6744; // @[icache.scala 135:42]
  wire [184:0] _GEN_10841 = replace & io_inst_sram_data_ok ? _GEN_9817 : _GEN_6745; // @[icache.scala 135:42]
  wire [184:0] _GEN_10842 = replace & io_inst_sram_data_ok ? _GEN_9818 : _GEN_6746; // @[icache.scala 135:42]
  wire [184:0] _GEN_10843 = replace & io_inst_sram_data_ok ? _GEN_9819 : _GEN_6747; // @[icache.scala 135:42]
  wire [184:0] _GEN_10844 = replace & io_inst_sram_data_ok ? _GEN_9820 : _GEN_6748; // @[icache.scala 135:42]
  wire [184:0] _GEN_10845 = replace & io_inst_sram_data_ok ? _GEN_9821 : _GEN_6749; // @[icache.scala 135:42]
  wire [184:0] _GEN_10846 = replace & io_inst_sram_data_ok ? _GEN_9822 : _GEN_6750; // @[icache.scala 135:42]
  wire [184:0] _GEN_10847 = replace & io_inst_sram_data_ok ? _GEN_9823 : _GEN_6751; // @[icache.scala 135:42]
  wire [184:0] _GEN_10848 = replace & io_inst_sram_data_ok ? _GEN_9824 : _GEN_6752; // @[icache.scala 135:42]
  wire [184:0] _GEN_10849 = replace & io_inst_sram_data_ok ? _GEN_9825 : _GEN_6753; // @[icache.scala 135:42]
  wire [184:0] _GEN_10850 = replace & io_inst_sram_data_ok ? _GEN_9826 : _GEN_6754; // @[icache.scala 135:42]
  wire [184:0] _GEN_10851 = replace & io_inst_sram_data_ok ? _GEN_9827 : _GEN_6755; // @[icache.scala 135:42]
  wire [184:0] _GEN_10852 = replace & io_inst_sram_data_ok ? _GEN_9828 : _GEN_6756; // @[icache.scala 135:42]
  wire [184:0] _GEN_10853 = replace & io_inst_sram_data_ok ? _GEN_9829 : _GEN_6757; // @[icache.scala 135:42]
  wire [184:0] _GEN_10854 = replace & io_inst_sram_data_ok ? _GEN_9830 : _GEN_6758; // @[icache.scala 135:42]
  wire [184:0] _GEN_10855 = replace & io_inst_sram_data_ok ? _GEN_9831 : _GEN_6759; // @[icache.scala 135:42]
  wire [184:0] _GEN_10856 = replace & io_inst_sram_data_ok ? _GEN_9832 : _GEN_6760; // @[icache.scala 135:42]
  wire [184:0] _GEN_10857 = replace & io_inst_sram_data_ok ? _GEN_9833 : _GEN_6761; // @[icache.scala 135:42]
  wire [184:0] _GEN_10858 = replace & io_inst_sram_data_ok ? _GEN_9834 : _GEN_6762; // @[icache.scala 135:42]
  wire [184:0] _GEN_10859 = replace & io_inst_sram_data_ok ? _GEN_9835 : _GEN_6763; // @[icache.scala 135:42]
  wire [184:0] _GEN_10860 = replace & io_inst_sram_data_ok ? _GEN_9836 : _GEN_6764; // @[icache.scala 135:42]
  wire [184:0] _GEN_10861 = replace & io_inst_sram_data_ok ? _GEN_9837 : _GEN_6765; // @[icache.scala 135:42]
  wire [184:0] _GEN_10862 = replace & io_inst_sram_data_ok ? _GEN_9838 : _GEN_6766; // @[icache.scala 135:42]
  wire [184:0] _GEN_10863 = replace & io_inst_sram_data_ok ? _GEN_9839 : _GEN_6767; // @[icache.scala 135:42]
  wire [184:0] _GEN_10864 = replace & io_inst_sram_data_ok ? _GEN_9840 : _GEN_6768; // @[icache.scala 135:42]
  wire [184:0] _GEN_10865 = replace & io_inst_sram_data_ok ? _GEN_9841 : _GEN_6769; // @[icache.scala 135:42]
  wire [184:0] _GEN_10866 = replace & io_inst_sram_data_ok ? _GEN_9842 : _GEN_6770; // @[icache.scala 135:42]
  wire [184:0] _GEN_10867 = replace & io_inst_sram_data_ok ? _GEN_9843 : _GEN_6771; // @[icache.scala 135:42]
  wire [184:0] _GEN_10868 = replace & io_inst_sram_data_ok ? _GEN_9844 : _GEN_6772; // @[icache.scala 135:42]
  wire [184:0] _GEN_10869 = replace & io_inst_sram_data_ok ? _GEN_9845 : _GEN_6773; // @[icache.scala 135:42]
  wire [184:0] _GEN_10870 = replace & io_inst_sram_data_ok ? _GEN_9846 : _GEN_6774; // @[icache.scala 135:42]
  wire [184:0] _GEN_10871 = replace & io_inst_sram_data_ok ? _GEN_9847 : _GEN_6775; // @[icache.scala 135:42]
  wire [184:0] _GEN_10872 = replace & io_inst_sram_data_ok ? _GEN_9848 : _GEN_6776; // @[icache.scala 135:42]
  wire [184:0] _GEN_10873 = replace & io_inst_sram_data_ok ? _GEN_9849 : _GEN_6777; // @[icache.scala 135:42]
  wire [184:0] _GEN_10874 = replace & io_inst_sram_data_ok ? _GEN_9850 : _GEN_6778; // @[icache.scala 135:42]
  wire [184:0] _GEN_10875 = replace & io_inst_sram_data_ok ? _GEN_9851 : _GEN_6779; // @[icache.scala 135:42]
  wire [184:0] _GEN_10876 = replace & io_inst_sram_data_ok ? _GEN_9852 : _GEN_6780; // @[icache.scala 135:42]
  wire [184:0] _GEN_10877 = replace & io_inst_sram_data_ok ? _GEN_9853 : _GEN_6781; // @[icache.scala 135:42]
  wire [184:0] _GEN_10878 = replace & io_inst_sram_data_ok ? _GEN_9854 : _GEN_6782; // @[icache.scala 135:42]
  wire [184:0] _GEN_10879 = replace & io_inst_sram_data_ok ? _GEN_9855 : _GEN_6783; // @[icache.scala 135:42]
  wire [184:0] _GEN_10880 = replace & io_inst_sram_data_ok ? _GEN_9856 : _GEN_6784; // @[icache.scala 135:42]
  wire [184:0] _GEN_10881 = replace & io_inst_sram_data_ok ? _GEN_9857 : _GEN_6785; // @[icache.scala 135:42]
  wire [184:0] _GEN_10882 = replace & io_inst_sram_data_ok ? _GEN_9858 : _GEN_6786; // @[icache.scala 135:42]
  wire [184:0] _GEN_10883 = replace & io_inst_sram_data_ok ? _GEN_9859 : _GEN_6787; // @[icache.scala 135:42]
  wire [184:0] _GEN_10884 = replace & io_inst_sram_data_ok ? _GEN_9860 : _GEN_6788; // @[icache.scala 135:42]
  wire [184:0] _GEN_10885 = replace & io_inst_sram_data_ok ? _GEN_9861 : _GEN_6789; // @[icache.scala 135:42]
  wire [184:0] _GEN_10886 = replace & io_inst_sram_data_ok ? _GEN_9862 : _GEN_6790; // @[icache.scala 135:42]
  wire [184:0] _GEN_10887 = replace & io_inst_sram_data_ok ? _GEN_9863 : _GEN_6791; // @[icache.scala 135:42]
  wire [184:0] _GEN_10888 = replace & io_inst_sram_data_ok ? _GEN_9864 : _GEN_6792; // @[icache.scala 135:42]
  wire [184:0] _GEN_10889 = replace & io_inst_sram_data_ok ? _GEN_9865 : _GEN_6793; // @[icache.scala 135:42]
  wire [184:0] _GEN_10890 = replace & io_inst_sram_data_ok ? _GEN_9866 : _GEN_6794; // @[icache.scala 135:42]
  wire [184:0] _GEN_10891 = replace & io_inst_sram_data_ok ? _GEN_9867 : _GEN_6795; // @[icache.scala 135:42]
  wire [184:0] _GEN_10892 = replace & io_inst_sram_data_ok ? _GEN_9868 : _GEN_6796; // @[icache.scala 135:42]
  wire [184:0] _GEN_10893 = replace & io_inst_sram_data_ok ? _GEN_9869 : _GEN_6797; // @[icache.scala 135:42]
  wire [184:0] _GEN_10894 = replace & io_inst_sram_data_ok ? _GEN_9870 : _GEN_6798; // @[icache.scala 135:42]
  wire [184:0] _GEN_10895 = replace & io_inst_sram_data_ok ? _GEN_9871 : _GEN_6799; // @[icache.scala 135:42]
  wire [184:0] _GEN_10896 = replace & io_inst_sram_data_ok ? _GEN_9872 : _GEN_6800; // @[icache.scala 135:42]
  wire [184:0] _GEN_10897 = replace & io_inst_sram_data_ok ? _GEN_9873 : _GEN_6801; // @[icache.scala 135:42]
  wire [184:0] _GEN_10898 = replace & io_inst_sram_data_ok ? _GEN_9874 : _GEN_6802; // @[icache.scala 135:42]
  wire [184:0] _GEN_10899 = replace & io_inst_sram_data_ok ? _GEN_9875 : _GEN_6803; // @[icache.scala 135:42]
  wire [184:0] _GEN_10900 = replace & io_inst_sram_data_ok ? _GEN_9876 : _GEN_6804; // @[icache.scala 135:42]
  wire [184:0] _GEN_10901 = replace & io_inst_sram_data_ok ? _GEN_9877 : _GEN_6805; // @[icache.scala 135:42]
  wire [184:0] _GEN_10902 = replace & io_inst_sram_data_ok ? _GEN_9878 : _GEN_6806; // @[icache.scala 135:42]
  wire [184:0] _GEN_10903 = replace & io_inst_sram_data_ok ? _GEN_9879 : _GEN_6807; // @[icache.scala 135:42]
  wire [184:0] _GEN_10904 = replace & io_inst_sram_data_ok ? _GEN_9880 : _GEN_6808; // @[icache.scala 135:42]
  wire [184:0] _GEN_10905 = replace & io_inst_sram_data_ok ? _GEN_9881 : _GEN_6809; // @[icache.scala 135:42]
  wire [184:0] _GEN_10906 = replace & io_inst_sram_data_ok ? _GEN_9882 : _GEN_6810; // @[icache.scala 135:42]
  wire [184:0] _GEN_10907 = replace & io_inst_sram_data_ok ? _GEN_9883 : _GEN_6811; // @[icache.scala 135:42]
  wire [184:0] _GEN_10908 = replace & io_inst_sram_data_ok ? _GEN_9884 : _GEN_6812; // @[icache.scala 135:42]
  wire [184:0] _GEN_10909 = replace & io_inst_sram_data_ok ? _GEN_9885 : _GEN_6813; // @[icache.scala 135:42]
  wire [184:0] _GEN_10910 = replace & io_inst_sram_data_ok ? _GEN_9886 : _GEN_6814; // @[icache.scala 135:42]
  wire [184:0] _GEN_10911 = replace & io_inst_sram_data_ok ? _GEN_9887 : _GEN_6815; // @[icache.scala 135:42]
  wire [184:0] _GEN_10912 = replace & io_inst_sram_data_ok ? _GEN_9888 : _GEN_6816; // @[icache.scala 135:42]
  wire [184:0] _GEN_10913 = replace & io_inst_sram_data_ok ? _GEN_9889 : _GEN_6817; // @[icache.scala 135:42]
  wire [184:0] _GEN_10914 = replace & io_inst_sram_data_ok ? _GEN_9890 : _GEN_6818; // @[icache.scala 135:42]
  wire [184:0] _GEN_10915 = replace & io_inst_sram_data_ok ? _GEN_9891 : _GEN_6819; // @[icache.scala 135:42]
  wire [184:0] _GEN_10916 = replace & io_inst_sram_data_ok ? _GEN_9892 : _GEN_6820; // @[icache.scala 135:42]
  wire [184:0] _GEN_10917 = replace & io_inst_sram_data_ok ? _GEN_9893 : _GEN_6821; // @[icache.scala 135:42]
  wire [184:0] _GEN_10918 = replace & io_inst_sram_data_ok ? _GEN_9894 : _GEN_6822; // @[icache.scala 135:42]
  wire [184:0] _GEN_10919 = replace & io_inst_sram_data_ok ? _GEN_9895 : _GEN_6823; // @[icache.scala 135:42]
  wire [184:0] _GEN_10920 = replace & io_inst_sram_data_ok ? _GEN_9896 : _GEN_6824; // @[icache.scala 135:42]
  wire [184:0] _GEN_10921 = replace & io_inst_sram_data_ok ? _GEN_9897 : _GEN_6825; // @[icache.scala 135:42]
  wire [184:0] _GEN_10922 = replace & io_inst_sram_data_ok ? _GEN_9898 : _GEN_6826; // @[icache.scala 135:42]
  wire [184:0] _GEN_10923 = replace & io_inst_sram_data_ok ? _GEN_9899 : _GEN_6827; // @[icache.scala 135:42]
  wire [184:0] _GEN_10924 = replace & io_inst_sram_data_ok ? _GEN_9900 : _GEN_6828; // @[icache.scala 135:42]
  wire [184:0] _GEN_10925 = replace & io_inst_sram_data_ok ? _GEN_9901 : _GEN_6829; // @[icache.scala 135:42]
  wire [184:0] _GEN_10926 = replace & io_inst_sram_data_ok ? _GEN_9902 : _GEN_6830; // @[icache.scala 135:42]
  wire [184:0] _GEN_10927 = replace & io_inst_sram_data_ok ? _GEN_9903 : _GEN_6831; // @[icache.scala 135:42]
  wire [184:0] _GEN_10928 = replace & io_inst_sram_data_ok ? _GEN_9904 : _GEN_6832; // @[icache.scala 135:42]
  wire [184:0] _GEN_10929 = replace & io_inst_sram_data_ok ? _GEN_9905 : _GEN_6833; // @[icache.scala 135:42]
  wire [184:0] _GEN_10930 = replace & io_inst_sram_data_ok ? _GEN_9906 : _GEN_6834; // @[icache.scala 135:42]
  wire [184:0] _GEN_10931 = replace & io_inst_sram_data_ok ? _GEN_9907 : _GEN_6835; // @[icache.scala 135:42]
  wire [184:0] _GEN_10932 = replace & io_inst_sram_data_ok ? _GEN_9908 : _GEN_6836; // @[icache.scala 135:42]
  wire [184:0] _GEN_10933 = replace & io_inst_sram_data_ok ? _GEN_9909 : _GEN_6837; // @[icache.scala 135:42]
  wire [184:0] _GEN_10934 = replace & io_inst_sram_data_ok ? _GEN_9910 : _GEN_6838; // @[icache.scala 135:42]
  wire [184:0] _GEN_10935 = replace & io_inst_sram_data_ok ? _GEN_9911 : _GEN_6839; // @[icache.scala 135:42]
  wire [184:0] _GEN_10936 = replace & io_inst_sram_data_ok ? _GEN_9912 : _GEN_6840; // @[icache.scala 135:42]
  wire [184:0] _GEN_10937 = replace & io_inst_sram_data_ok ? _GEN_9913 : _GEN_6841; // @[icache.scala 135:42]
  wire [184:0] _GEN_10938 = replace & io_inst_sram_data_ok ? _GEN_9914 : _GEN_6842; // @[icache.scala 135:42]
  wire [184:0] _GEN_10939 = replace & io_inst_sram_data_ok ? _GEN_9915 : _GEN_6843; // @[icache.scala 135:42]
  wire [184:0] _GEN_10940 = replace & io_inst_sram_data_ok ? _GEN_9916 : _GEN_6844; // @[icache.scala 135:42]
  wire [184:0] _GEN_10941 = replace & io_inst_sram_data_ok ? _GEN_9917 : _GEN_6845; // @[icache.scala 135:42]
  wire [184:0] _GEN_10942 = replace & io_inst_sram_data_ok ? _GEN_9918 : _GEN_6846; // @[icache.scala 135:42]
  wire [184:0] _GEN_10943 = replace & io_inst_sram_data_ok ? _GEN_9919 : _GEN_6847; // @[icache.scala 135:42]
  wire [184:0] _GEN_10944 = replace & io_inst_sram_data_ok ? _GEN_9920 : _GEN_6848; // @[icache.scala 135:42]
  wire [184:0] _GEN_10945 = replace & io_inst_sram_data_ok ? _GEN_9921 : _GEN_6849; // @[icache.scala 135:42]
  wire [184:0] _GEN_10946 = replace & io_inst_sram_data_ok ? _GEN_9922 : _GEN_6850; // @[icache.scala 135:42]
  wire [184:0] _GEN_10947 = replace & io_inst_sram_data_ok ? _GEN_9923 : _GEN_6851; // @[icache.scala 135:42]
  wire [184:0] _GEN_10948 = replace & io_inst_sram_data_ok ? _GEN_9924 : _GEN_6852; // @[icache.scala 135:42]
  wire [184:0] _GEN_10949 = replace & io_inst_sram_data_ok ? _GEN_9925 : _GEN_6853; // @[icache.scala 135:42]
  wire [184:0] _GEN_10950 = replace & io_inst_sram_data_ok ? _GEN_9926 : _GEN_6854; // @[icache.scala 135:42]
  wire [184:0] _GEN_10951 = replace & io_inst_sram_data_ok ? _GEN_9927 : _GEN_6855; // @[icache.scala 135:42]
  wire [184:0] _GEN_10952 = replace & io_inst_sram_data_ok ? _GEN_9928 : _GEN_6856; // @[icache.scala 135:42]
  wire [184:0] _GEN_10953 = replace & io_inst_sram_data_ok ? _GEN_9929 : _GEN_6857; // @[icache.scala 135:42]
  wire [184:0] _GEN_10954 = replace & io_inst_sram_data_ok ? _GEN_9930 : _GEN_6858; // @[icache.scala 135:42]
  wire [184:0] _GEN_10955 = replace & io_inst_sram_data_ok ? _GEN_9931 : _GEN_6859; // @[icache.scala 135:42]
  wire [184:0] _GEN_10956 = replace & io_inst_sram_data_ok ? _GEN_9932 : _GEN_6860; // @[icache.scala 135:42]
  wire [184:0] _GEN_10957 = replace & io_inst_sram_data_ok ? _GEN_9933 : _GEN_6861; // @[icache.scala 135:42]
  wire [184:0] _GEN_10958 = replace & io_inst_sram_data_ok ? _GEN_9934 : _GEN_6862; // @[icache.scala 135:42]
  wire [184:0] _GEN_10959 = replace & io_inst_sram_data_ok ? _GEN_9935 : _GEN_6863; // @[icache.scala 135:42]
  wire [184:0] _GEN_10960 = replace & io_inst_sram_data_ok ? _GEN_9936 : _GEN_6864; // @[icache.scala 135:42]
  wire [184:0] _GEN_10961 = replace & io_inst_sram_data_ok ? _GEN_9937 : _GEN_6865; // @[icache.scala 135:42]
  wire [184:0] _GEN_10962 = replace & io_inst_sram_data_ok ? _GEN_9938 : _GEN_6866; // @[icache.scala 135:42]
  wire [184:0] _GEN_10963 = replace & io_inst_sram_data_ok ? _GEN_9939 : _GEN_6867; // @[icache.scala 135:42]
  wire [184:0] _GEN_10964 = replace & io_inst_sram_data_ok ? _GEN_9940 : _GEN_6868; // @[icache.scala 135:42]
  wire [184:0] _GEN_10965 = replace & io_inst_sram_data_ok ? _GEN_9941 : _GEN_6869; // @[icache.scala 135:42]
  wire [184:0] _GEN_10966 = replace & io_inst_sram_data_ok ? _GEN_9942 : _GEN_6870; // @[icache.scala 135:42]
  wire [184:0] _GEN_10967 = replace & io_inst_sram_data_ok ? _GEN_9943 : _GEN_6871; // @[icache.scala 135:42]
  wire [184:0] _GEN_10968 = replace & io_inst_sram_data_ok ? _GEN_9944 : _GEN_6872; // @[icache.scala 135:42]
  wire [184:0] _GEN_10969 = replace & io_inst_sram_data_ok ? _GEN_9945 : _GEN_6873; // @[icache.scala 135:42]
  wire [184:0] _GEN_10970 = replace & io_inst_sram_data_ok ? _GEN_9946 : _GEN_6874; // @[icache.scala 135:42]
  wire [184:0] _GEN_10971 = replace & io_inst_sram_data_ok ? _GEN_9947 : _GEN_6875; // @[icache.scala 135:42]
  wire [184:0] _GEN_10972 = replace & io_inst_sram_data_ok ? _GEN_9948 : _GEN_6876; // @[icache.scala 135:42]
  wire [184:0] _GEN_10973 = replace & io_inst_sram_data_ok ? _GEN_9949 : _GEN_6877; // @[icache.scala 135:42]
  wire [184:0] _GEN_10974 = replace & io_inst_sram_data_ok ? _GEN_9950 : _GEN_6878; // @[icache.scala 135:42]
  wire [184:0] _GEN_10975 = replace & io_inst_sram_data_ok ? _GEN_9951 : _GEN_6879; // @[icache.scala 135:42]
  wire [184:0] _GEN_10976 = replace & io_inst_sram_data_ok ? _GEN_9952 : _GEN_6880; // @[icache.scala 135:42]
  wire [184:0] _GEN_10977 = replace & io_inst_sram_data_ok ? _GEN_9953 : _GEN_6881; // @[icache.scala 135:42]
  wire [184:0] _GEN_10978 = replace & io_inst_sram_data_ok ? _GEN_9954 : _GEN_6882; // @[icache.scala 135:42]
  wire [184:0] _GEN_10979 = replace & io_inst_sram_data_ok ? _GEN_9955 : _GEN_6883; // @[icache.scala 135:42]
  wire [184:0] _GEN_10980 = replace & io_inst_sram_data_ok ? _GEN_9956 : _GEN_6884; // @[icache.scala 135:42]
  wire [184:0] _GEN_10981 = replace & io_inst_sram_data_ok ? _GEN_9957 : _GEN_6885; // @[icache.scala 135:42]
  wire [184:0] _GEN_10982 = replace & io_inst_sram_data_ok ? _GEN_9958 : _GEN_6886; // @[icache.scala 135:42]
  wire [184:0] _GEN_10983 = replace & io_inst_sram_data_ok ? _GEN_9959 : _GEN_6887; // @[icache.scala 135:42]
  wire [184:0] _GEN_10984 = replace & io_inst_sram_data_ok ? _GEN_9960 : _GEN_6888; // @[icache.scala 135:42]
  wire [184:0] _GEN_10985 = replace & io_inst_sram_data_ok ? _GEN_9961 : _GEN_6889; // @[icache.scala 135:42]
  wire [184:0] _GEN_10986 = replace & io_inst_sram_data_ok ? _GEN_9962 : _GEN_6890; // @[icache.scala 135:42]
  wire [184:0] _GEN_10987 = replace & io_inst_sram_data_ok ? _GEN_9963 : _GEN_6891; // @[icache.scala 135:42]
  wire [184:0] _GEN_10988 = replace & io_inst_sram_data_ok ? _GEN_9964 : _GEN_6892; // @[icache.scala 135:42]
  wire [184:0] _GEN_10989 = replace & io_inst_sram_data_ok ? _GEN_9965 : _GEN_6893; // @[icache.scala 135:42]
  wire [184:0] _GEN_10990 = replace & io_inst_sram_data_ok ? _GEN_9966 : _GEN_6894; // @[icache.scala 135:42]
  wire [184:0] _GEN_10991 = replace & io_inst_sram_data_ok ? _GEN_9967 : _GEN_6895; // @[icache.scala 135:42]
  wire [184:0] _GEN_10992 = replace & io_inst_sram_data_ok ? _GEN_9968 : _GEN_6896; // @[icache.scala 135:42]
  wire [184:0] _GEN_10993 = replace & io_inst_sram_data_ok ? _GEN_9969 : _GEN_6897; // @[icache.scala 135:42]
  wire [184:0] _GEN_10994 = replace & io_inst_sram_data_ok ? _GEN_9970 : _GEN_6898; // @[icache.scala 135:42]
  wire [184:0] _GEN_10995 = replace & io_inst_sram_data_ok ? _GEN_9971 : _GEN_6899; // @[icache.scala 135:42]
  wire [184:0] _GEN_10996 = replace & io_inst_sram_data_ok ? _GEN_9972 : _GEN_6900; // @[icache.scala 135:42]
  wire [184:0] _GEN_10997 = replace & io_inst_sram_data_ok ? _GEN_9973 : _GEN_6901; // @[icache.scala 135:42]
  wire [184:0] _GEN_10998 = replace & io_inst_sram_data_ok ? _GEN_9974 : _GEN_6902; // @[icache.scala 135:42]
  wire [184:0] _GEN_10999 = replace & io_inst_sram_data_ok ? _GEN_9975 : _GEN_6903; // @[icache.scala 135:42]
  wire [184:0] _GEN_11000 = replace & io_inst_sram_data_ok ? _GEN_9976 : _GEN_6904; // @[icache.scala 135:42]
  wire [184:0] _GEN_11001 = replace & io_inst_sram_data_ok ? _GEN_9977 : _GEN_6905; // @[icache.scala 135:42]
  wire [184:0] _GEN_11002 = replace & io_inst_sram_data_ok ? _GEN_9978 : _GEN_6906; // @[icache.scala 135:42]
  wire [184:0] _GEN_11003 = replace & io_inst_sram_data_ok ? _GEN_9979 : _GEN_6907; // @[icache.scala 135:42]
  wire [184:0] _GEN_11004 = replace & io_inst_sram_data_ok ? _GEN_9980 : _GEN_6908; // @[icache.scala 135:42]
  wire [184:0] _GEN_11005 = replace & io_inst_sram_data_ok ? _GEN_9981 : _GEN_6909; // @[icache.scala 135:42]
  wire [184:0] _GEN_11006 = replace & io_inst_sram_data_ok ? _GEN_9982 : _GEN_6910; // @[icache.scala 135:42]
  wire [184:0] _GEN_11007 = replace & io_inst_sram_data_ok ? _GEN_9983 : _GEN_6911; // @[icache.scala 135:42]
  wire [184:0] _GEN_11008 = replace & io_inst_sram_data_ok ? _GEN_9984 : _GEN_6912; // @[icache.scala 135:42]
  wire [184:0] _GEN_11009 = replace & io_inst_sram_data_ok ? _GEN_9985 : _GEN_6913; // @[icache.scala 135:42]
  wire [184:0] _GEN_11010 = replace & io_inst_sram_data_ok ? _GEN_9986 : _GEN_6914; // @[icache.scala 135:42]
  wire [184:0] _GEN_11011 = replace & io_inst_sram_data_ok ? _GEN_9987 : _GEN_6915; // @[icache.scala 135:42]
  wire [184:0] _GEN_11012 = replace & io_inst_sram_data_ok ? _GEN_9988 : _GEN_6916; // @[icache.scala 135:42]
  wire [184:0] _GEN_11013 = replace & io_inst_sram_data_ok ? _GEN_9989 : _GEN_6917; // @[icache.scala 135:42]
  wire [184:0] _GEN_11014 = replace & io_inst_sram_data_ok ? _GEN_9990 : _GEN_6918; // @[icache.scala 135:42]
  wire [184:0] _GEN_11015 = replace & io_inst_sram_data_ok ? _GEN_9991 : _GEN_6919; // @[icache.scala 135:42]
  wire [184:0] _GEN_11016 = replace & io_inst_sram_data_ok ? _GEN_9992 : _GEN_6920; // @[icache.scala 135:42]
  wire [184:0] _GEN_11017 = replace & io_inst_sram_data_ok ? _GEN_9993 : _GEN_6921; // @[icache.scala 135:42]
  wire [184:0] _GEN_11018 = replace & io_inst_sram_data_ok ? _GEN_9994 : _GEN_6922; // @[icache.scala 135:42]
  wire [184:0] _GEN_11019 = replace & io_inst_sram_data_ok ? _GEN_9995 : _GEN_6923; // @[icache.scala 135:42]
  wire [184:0] _GEN_11020 = replace & io_inst_sram_data_ok ? _GEN_9996 : _GEN_6924; // @[icache.scala 135:42]
  wire [184:0] _GEN_11021 = replace & io_inst_sram_data_ok ? _GEN_9997 : _GEN_6925; // @[icache.scala 135:42]
  wire [184:0] _GEN_11022 = replace & io_inst_sram_data_ok ? _GEN_9998 : _GEN_6926; // @[icache.scala 135:42]
  wire [184:0] _GEN_11023 = replace & io_inst_sram_data_ok ? _GEN_9999 : _GEN_6927; // @[icache.scala 135:42]
  wire [184:0] _GEN_11024 = replace & io_inst_sram_data_ok ? _GEN_10000 : _GEN_6928; // @[icache.scala 135:42]
  wire [184:0] _GEN_11025 = replace & io_inst_sram_data_ok ? _GEN_10001 : _GEN_6929; // @[icache.scala 135:42]
  wire [184:0] _GEN_11026 = replace & io_inst_sram_data_ok ? _GEN_10002 : _GEN_6930; // @[icache.scala 135:42]
  wire [184:0] _GEN_11027 = replace & io_inst_sram_data_ok ? _GEN_10003 : _GEN_6931; // @[icache.scala 135:42]
  wire [184:0] _GEN_11028 = replace & io_inst_sram_data_ok ? _GEN_10004 : _GEN_6932; // @[icache.scala 135:42]
  wire [184:0] _GEN_11029 = replace & io_inst_sram_data_ok ? _GEN_10005 : _GEN_6933; // @[icache.scala 135:42]
  wire [184:0] _GEN_11030 = replace & io_inst_sram_data_ok ? _GEN_10006 : _GEN_6934; // @[icache.scala 135:42]
  wire [184:0] _GEN_11031 = replace & io_inst_sram_data_ok ? _GEN_10007 : _GEN_6935; // @[icache.scala 135:42]
  wire [184:0] _GEN_11032 = replace & io_inst_sram_data_ok ? _GEN_10008 : _GEN_6936; // @[icache.scala 135:42]
  wire [184:0] _GEN_11033 = replace & io_inst_sram_data_ok ? _GEN_10009 : _GEN_6937; // @[icache.scala 135:42]
  wire [184:0] _GEN_11034 = replace & io_inst_sram_data_ok ? _GEN_10010 : _GEN_6938; // @[icache.scala 135:42]
  wire [184:0] _GEN_11035 = replace & io_inst_sram_data_ok ? _GEN_10011 : _GEN_6939; // @[icache.scala 135:42]
  wire [184:0] _GEN_11036 = replace & io_inst_sram_data_ok ? _GEN_10012 : _GEN_6940; // @[icache.scala 135:42]
  wire [184:0] _GEN_11037 = replace & io_inst_sram_data_ok ? _GEN_10013 : _GEN_6941; // @[icache.scala 135:42]
  wire [184:0] _GEN_11038 = replace & io_inst_sram_data_ok ? _GEN_10014 : _GEN_6942; // @[icache.scala 135:42]
  wire [184:0] _GEN_11039 = replace & io_inst_sram_data_ok ? _GEN_10015 : _GEN_6943; // @[icache.scala 135:42]
  wire [184:0] _GEN_11040 = replace & io_inst_sram_data_ok ? _GEN_10016 : _GEN_6944; // @[icache.scala 135:42]
  wire [184:0] _GEN_11041 = replace & io_inst_sram_data_ok ? _GEN_10017 : _GEN_6945; // @[icache.scala 135:42]
  wire [184:0] _GEN_11042 = replace & io_inst_sram_data_ok ? _GEN_10018 : _GEN_6946; // @[icache.scala 135:42]
  wire [184:0] _GEN_11043 = replace & io_inst_sram_data_ok ? _GEN_10019 : _GEN_6947; // @[icache.scala 135:42]
  wire [184:0] _GEN_11044 = replace & io_inst_sram_data_ok ? _GEN_10020 : _GEN_6948; // @[icache.scala 135:42]
  wire [184:0] _GEN_11045 = replace & io_inst_sram_data_ok ? _GEN_10021 : _GEN_6949; // @[icache.scala 135:42]
  wire [184:0] _GEN_11046 = replace & io_inst_sram_data_ok ? _GEN_10022 : _GEN_6950; // @[icache.scala 135:42]
  wire [184:0] _GEN_11047 = replace & io_inst_sram_data_ok ? _GEN_10023 : _GEN_6951; // @[icache.scala 135:42]
  wire [184:0] _GEN_11048 = replace & io_inst_sram_data_ok ? _GEN_10024 : _GEN_6952; // @[icache.scala 135:42]
  wire [184:0] _GEN_11049 = replace & io_inst_sram_data_ok ? _GEN_10025 : _GEN_6953; // @[icache.scala 135:42]
  wire [184:0] _GEN_11050 = replace & io_inst_sram_data_ok ? _GEN_10026 : _GEN_6954; // @[icache.scala 135:42]
  wire [184:0] _GEN_11051 = replace & io_inst_sram_data_ok ? _GEN_10027 : _GEN_6955; // @[icache.scala 135:42]
  wire [184:0] _GEN_11052 = replace & io_inst_sram_data_ok ? _GEN_10028 : _GEN_6956; // @[icache.scala 135:42]
  wire [184:0] _GEN_11053 = replace & io_inst_sram_data_ok ? _GEN_10029 : _GEN_6957; // @[icache.scala 135:42]
  wire [184:0] _GEN_11054 = replace & io_inst_sram_data_ok ? _GEN_10030 : _GEN_6958; // @[icache.scala 135:42]
  wire [184:0] _GEN_11055 = replace & io_inst_sram_data_ok ? _GEN_10031 : _GEN_6959; // @[icache.scala 135:42]
  wire [184:0] _GEN_11056 = replace & io_inst_sram_data_ok ? _GEN_10032 : _GEN_6960; // @[icache.scala 135:42]
  wire [184:0] _GEN_11057 = replace & io_inst_sram_data_ok ? _GEN_10033 : _GEN_6961; // @[icache.scala 135:42]
  wire [184:0] _GEN_11058 = replace & io_inst_sram_data_ok ? _GEN_10034 : _GEN_6962; // @[icache.scala 135:42]
  wire [184:0] _GEN_11059 = replace & io_inst_sram_data_ok ? _GEN_10035 : _GEN_6963; // @[icache.scala 135:42]
  wire [184:0] _GEN_11060 = replace & io_inst_sram_data_ok ? _GEN_10036 : _GEN_6964; // @[icache.scala 135:42]
  wire [184:0] _GEN_11061 = replace & io_inst_sram_data_ok ? _GEN_10037 : _GEN_6965; // @[icache.scala 135:42]
  wire [184:0] _GEN_11062 = replace & io_inst_sram_data_ok ? _GEN_10038 : _GEN_6966; // @[icache.scala 135:42]
  wire [184:0] _GEN_11063 = replace & io_inst_sram_data_ok ? _GEN_10039 : _GEN_6967; // @[icache.scala 135:42]
  wire [184:0] _GEN_11064 = replace & io_inst_sram_data_ok ? _GEN_10040 : _GEN_6968; // @[icache.scala 135:42]
  wire [184:0] _GEN_11065 = replace & io_inst_sram_data_ok ? _GEN_10041 : _GEN_6969; // @[icache.scala 135:42]
  wire [184:0] _GEN_11066 = replace & io_inst_sram_data_ok ? _GEN_10042 : _GEN_6970; // @[icache.scala 135:42]
  wire [184:0] _GEN_11067 = replace & io_inst_sram_data_ok ? _GEN_10043 : _GEN_6971; // @[icache.scala 135:42]
  wire [184:0] _GEN_11068 = replace & io_inst_sram_data_ok ? _GEN_10044 : _GEN_6972; // @[icache.scala 135:42]
  wire [184:0] _GEN_11069 = replace & io_inst_sram_data_ok ? _GEN_10045 : _GEN_6973; // @[icache.scala 135:42]
  wire [184:0] _GEN_11070 = replace & io_inst_sram_data_ok ? _GEN_10046 : _GEN_6974; // @[icache.scala 135:42]
  wire [184:0] _GEN_11071 = replace & io_inst_sram_data_ok ? _GEN_10047 : _GEN_6975; // @[icache.scala 135:42]
  wire [184:0] _GEN_11072 = replace & io_inst_sram_data_ok ? _GEN_10048 : _GEN_6976; // @[icache.scala 135:42]
  wire [184:0] _GEN_11073 = replace & io_inst_sram_data_ok ? _GEN_10049 : _GEN_6977; // @[icache.scala 135:42]
  wire [184:0] _GEN_11074 = replace & io_inst_sram_data_ok ? _GEN_10050 : _GEN_6978; // @[icache.scala 135:42]
  wire [184:0] _GEN_11075 = replace & io_inst_sram_data_ok ? _GEN_10051 : _GEN_6979; // @[icache.scala 135:42]
  wire [184:0] _GEN_11076 = replace & io_inst_sram_data_ok ? _GEN_10052 : _GEN_6980; // @[icache.scala 135:42]
  wire [184:0] _GEN_11077 = replace & io_inst_sram_data_ok ? _GEN_10053 : _GEN_6981; // @[icache.scala 135:42]
  wire [184:0] _GEN_11078 = replace & io_inst_sram_data_ok ? _GEN_10054 : _GEN_6982; // @[icache.scala 135:42]
  wire [184:0] _GEN_11079 = replace & io_inst_sram_data_ok ? _GEN_10055 : _GEN_6983; // @[icache.scala 135:42]
  wire [184:0] _GEN_11080 = replace & io_inst_sram_data_ok ? _GEN_10056 : _GEN_6984; // @[icache.scala 135:42]
  wire [184:0] _GEN_11081 = replace & io_inst_sram_data_ok ? _GEN_10057 : _GEN_6985; // @[icache.scala 135:42]
  wire [184:0] _GEN_11082 = replace & io_inst_sram_data_ok ? _GEN_10058 : _GEN_6986; // @[icache.scala 135:42]
  wire [184:0] _GEN_11083 = replace & io_inst_sram_data_ok ? _GEN_10059 : _GEN_6987; // @[icache.scala 135:42]
  wire [184:0] _GEN_11084 = replace & io_inst_sram_data_ok ? _GEN_10060 : _GEN_6988; // @[icache.scala 135:42]
  wire [184:0] _GEN_11085 = replace & io_inst_sram_data_ok ? _GEN_10061 : _GEN_6989; // @[icache.scala 135:42]
  wire [184:0] _GEN_11086 = replace & io_inst_sram_data_ok ? _GEN_10062 : _GEN_6990; // @[icache.scala 135:42]
  wire [184:0] _GEN_11087 = replace & io_inst_sram_data_ok ? _GEN_10063 : _GEN_6991; // @[icache.scala 135:42]
  wire [184:0] _GEN_11088 = replace & io_inst_sram_data_ok ? _GEN_10064 : _GEN_6992; // @[icache.scala 135:42]
  wire [184:0] _GEN_11089 = replace & io_inst_sram_data_ok ? _GEN_10065 : _GEN_6993; // @[icache.scala 135:42]
  wire [184:0] _GEN_11090 = replace & io_inst_sram_data_ok ? _GEN_10066 : _GEN_6994; // @[icache.scala 135:42]
  wire [184:0] _GEN_11091 = replace & io_inst_sram_data_ok ? _GEN_10067 : _GEN_6995; // @[icache.scala 135:42]
  wire [184:0] _GEN_11092 = replace & io_inst_sram_data_ok ? _GEN_10068 : _GEN_6996; // @[icache.scala 135:42]
  wire [184:0] _GEN_11093 = replace & io_inst_sram_data_ok ? _GEN_10069 : _GEN_6997; // @[icache.scala 135:42]
  wire [184:0] _GEN_11094 = replace & io_inst_sram_data_ok ? _GEN_10070 : _GEN_6998; // @[icache.scala 135:42]
  wire [184:0] _GEN_11095 = replace & io_inst_sram_data_ok ? _GEN_10071 : _GEN_6999; // @[icache.scala 135:42]
  wire [184:0] _GEN_11096 = replace & io_inst_sram_data_ok ? _GEN_10072 : _GEN_7000; // @[icache.scala 135:42]
  wire [184:0] _GEN_11097 = replace & io_inst_sram_data_ok ? _GEN_10073 : _GEN_7001; // @[icache.scala 135:42]
  wire [184:0] _GEN_11098 = replace & io_inst_sram_data_ok ? _GEN_10074 : _GEN_7002; // @[icache.scala 135:42]
  wire [184:0] _GEN_11099 = replace & io_inst_sram_data_ok ? _GEN_10075 : _GEN_7003; // @[icache.scala 135:42]
  wire [184:0] _GEN_11100 = replace & io_inst_sram_data_ok ? _GEN_10076 : _GEN_7004; // @[icache.scala 135:42]
  wire [184:0] _GEN_11101 = replace & io_inst_sram_data_ok ? _GEN_10077 : _GEN_7005; // @[icache.scala 135:42]
  wire [184:0] _GEN_11102 = replace & io_inst_sram_data_ok ? _GEN_10078 : _GEN_7006; // @[icache.scala 135:42]
  wire [184:0] _GEN_11103 = replace & io_inst_sram_data_ok ? _GEN_10079 : _GEN_7007; // @[icache.scala 135:42]
  wire [184:0] _GEN_11104 = replace & io_inst_sram_data_ok ? _GEN_10080 : _GEN_7008; // @[icache.scala 135:42]
  wire [184:0] _GEN_11105 = replace & io_inst_sram_data_ok ? _GEN_10081 : _GEN_7009; // @[icache.scala 135:42]
  wire [184:0] _GEN_11106 = replace & io_inst_sram_data_ok ? _GEN_10082 : _GEN_7010; // @[icache.scala 135:42]
  wire [184:0] _GEN_11107 = replace & io_inst_sram_data_ok ? _GEN_10083 : _GEN_7011; // @[icache.scala 135:42]
  wire [184:0] _GEN_11108 = replace & io_inst_sram_data_ok ? _GEN_10084 : _GEN_7012; // @[icache.scala 135:42]
  wire [184:0] _GEN_11109 = replace & io_inst_sram_data_ok ? _GEN_10085 : _GEN_7013; // @[icache.scala 135:42]
  wire [184:0] _GEN_11110 = replace & io_inst_sram_data_ok ? _GEN_10086 : _GEN_7014; // @[icache.scala 135:42]
  wire [184:0] _GEN_11111 = replace & io_inst_sram_data_ok ? _GEN_10087 : _GEN_7015; // @[icache.scala 135:42]
  wire [184:0] _GEN_11112 = replace & io_inst_sram_data_ok ? _GEN_10088 : _GEN_7016; // @[icache.scala 135:42]
  wire [184:0] _GEN_11113 = replace & io_inst_sram_data_ok ? _GEN_10089 : _GEN_7017; // @[icache.scala 135:42]
  wire [184:0] _GEN_11114 = replace & io_inst_sram_data_ok ? _GEN_10090 : _GEN_7018; // @[icache.scala 135:42]
  wire [184:0] _GEN_11115 = replace & io_inst_sram_data_ok ? _GEN_10091 : _GEN_7019; // @[icache.scala 135:42]
  wire [184:0] _GEN_11116 = replace & io_inst_sram_data_ok ? _GEN_10092 : _GEN_7020; // @[icache.scala 135:42]
  wire [184:0] _GEN_11117 = replace & io_inst_sram_data_ok ? _GEN_10093 : _GEN_7021; // @[icache.scala 135:42]
  wire [184:0] _GEN_11118 = replace & io_inst_sram_data_ok ? _GEN_10094 : _GEN_7022; // @[icache.scala 135:42]
  wire [184:0] _GEN_11119 = replace & io_inst_sram_data_ok ? _GEN_10095 : _GEN_7023; // @[icache.scala 135:42]
  wire [184:0] _GEN_11120 = replace & io_inst_sram_data_ok ? _GEN_10096 : _GEN_7024; // @[icache.scala 135:42]
  wire [184:0] _GEN_11121 = replace & io_inst_sram_data_ok ? _GEN_10097 : _GEN_7025; // @[icache.scala 135:42]
  wire [184:0] _GEN_11122 = replace & io_inst_sram_data_ok ? _GEN_10098 : _GEN_7026; // @[icache.scala 135:42]
  wire [184:0] _GEN_11123 = replace & io_inst_sram_data_ok ? _GEN_10099 : _GEN_7027; // @[icache.scala 135:42]
  wire [184:0] _GEN_11124 = replace & io_inst_sram_data_ok ? _GEN_10100 : _GEN_7028; // @[icache.scala 135:42]
  wire [184:0] _GEN_11125 = replace & io_inst_sram_data_ok ? _GEN_10101 : _GEN_7029; // @[icache.scala 135:42]
  wire [184:0] _GEN_11126 = replace & io_inst_sram_data_ok ? _GEN_10102 : _GEN_7030; // @[icache.scala 135:42]
  wire [184:0] _GEN_11127 = replace & io_inst_sram_data_ok ? _GEN_10103 : _GEN_7031; // @[icache.scala 135:42]
  wire [184:0] _GEN_11128 = replace & io_inst_sram_data_ok ? _GEN_10104 : _GEN_7032; // @[icache.scala 135:42]
  wire [184:0] _GEN_11129 = replace & io_inst_sram_data_ok ? _GEN_10105 : _GEN_7033; // @[icache.scala 135:42]
  wire [184:0] _GEN_11130 = replace & io_inst_sram_data_ok ? _GEN_10106 : _GEN_7034; // @[icache.scala 135:42]
  wire [184:0] _GEN_11131 = replace & io_inst_sram_data_ok ? _GEN_10107 : _GEN_7035; // @[icache.scala 135:42]
  wire [184:0] _GEN_11132 = replace & io_inst_sram_data_ok ? _GEN_10108 : _GEN_7036; // @[icache.scala 135:42]
  wire [184:0] _GEN_11133 = replace & io_inst_sram_data_ok ? _GEN_10109 : _GEN_7037; // @[icache.scala 135:42]
  wire [184:0] _GEN_11134 = replace & io_inst_sram_data_ok ? _GEN_10110 : _GEN_7038; // @[icache.scala 135:42]
  wire [184:0] _GEN_11135 = replace & io_inst_sram_data_ok ? _GEN_10111 : _GEN_7039; // @[icache.scala 135:42]
  wire [184:0] _GEN_11136 = replace & io_inst_sram_data_ok ? _GEN_10112 : _GEN_7040; // @[icache.scala 135:42]
  wire [184:0] _GEN_11137 = replace & io_inst_sram_data_ok ? _GEN_10113 : _GEN_7041; // @[icache.scala 135:42]
  wire [184:0] _GEN_11138 = replace & io_inst_sram_data_ok ? _GEN_10114 : _GEN_7042; // @[icache.scala 135:42]
  wire [184:0] _GEN_11139 = replace & io_inst_sram_data_ok ? _GEN_10115 : _GEN_7043; // @[icache.scala 135:42]
  wire [184:0] _GEN_11140 = replace & io_inst_sram_data_ok ? _GEN_10116 : _GEN_7044; // @[icache.scala 135:42]
  wire [184:0] _GEN_11141 = replace & io_inst_sram_data_ok ? _GEN_10117 : _GEN_7045; // @[icache.scala 135:42]
  wire [184:0] _GEN_11142 = replace & io_inst_sram_data_ok ? _GEN_10118 : _GEN_7046; // @[icache.scala 135:42]
  wire [184:0] _GEN_11143 = replace & io_inst_sram_data_ok ? _GEN_10119 : _GEN_7047; // @[icache.scala 135:42]
  wire [184:0] _GEN_11144 = replace & io_inst_sram_data_ok ? _GEN_10120 : _GEN_7048; // @[icache.scala 135:42]
  wire [184:0] _GEN_11145 = replace & io_inst_sram_data_ok ? _GEN_10121 : _GEN_7049; // @[icache.scala 135:42]
  wire [184:0] _GEN_11146 = replace & io_inst_sram_data_ok ? _GEN_10122 : _GEN_7050; // @[icache.scala 135:42]
  wire [184:0] _GEN_11147 = replace & io_inst_sram_data_ok ? _GEN_10123 : _GEN_7051; // @[icache.scala 135:42]
  wire [184:0] _GEN_11148 = replace & io_inst_sram_data_ok ? _GEN_10124 : _GEN_7052; // @[icache.scala 135:42]
  wire [184:0] _GEN_11149 = replace & io_inst_sram_data_ok ? _GEN_10125 : _GEN_7053; // @[icache.scala 135:42]
  wire [184:0] _GEN_11150 = replace & io_inst_sram_data_ok ? _GEN_10126 : _GEN_7054; // @[icache.scala 135:42]
  wire [184:0] _GEN_11151 = replace & io_inst_sram_data_ok ? _GEN_10127 : _GEN_7055; // @[icache.scala 135:42]
  wire [184:0] _GEN_11152 = replace & io_inst_sram_data_ok ? _GEN_10128 : _GEN_7056; // @[icache.scala 135:42]
  wire [184:0] _GEN_11153 = replace & io_inst_sram_data_ok ? _GEN_10129 : _GEN_7057; // @[icache.scala 135:42]
  wire [184:0] _GEN_11154 = replace & io_inst_sram_data_ok ? _GEN_10130 : _GEN_7058; // @[icache.scala 135:42]
  wire [184:0] _GEN_11155 = replace & io_inst_sram_data_ok ? _GEN_10131 : _GEN_7059; // @[icache.scala 135:42]
  wire [184:0] _GEN_11156 = replace & io_inst_sram_data_ok ? _GEN_10132 : _GEN_7060; // @[icache.scala 135:42]
  wire [184:0] _GEN_11157 = replace & io_inst_sram_data_ok ? _GEN_10133 : _GEN_7061; // @[icache.scala 135:42]
  wire [184:0] _GEN_11158 = replace & io_inst_sram_data_ok ? _GEN_10134 : _GEN_7062; // @[icache.scala 135:42]
  wire [184:0] _GEN_11159 = replace & io_inst_sram_data_ok ? _GEN_10135 : _GEN_7063; // @[icache.scala 135:42]
  wire [184:0] _GEN_11160 = replace & io_inst_sram_data_ok ? _GEN_10136 : _GEN_7064; // @[icache.scala 135:42]
  wire [184:0] _GEN_11161 = replace & io_inst_sram_data_ok ? _GEN_10137 : _GEN_7065; // @[icache.scala 135:42]
  wire [184:0] _GEN_11162 = replace & io_inst_sram_data_ok ? _GEN_10138 : _GEN_7066; // @[icache.scala 135:42]
  wire [184:0] _GEN_11163 = replace & io_inst_sram_data_ok ? _GEN_10139 : _GEN_7067; // @[icache.scala 135:42]
  wire [184:0] _GEN_11164 = replace & io_inst_sram_data_ok ? _GEN_10140 : _GEN_7068; // @[icache.scala 135:42]
  wire [184:0] _GEN_11165 = replace & io_inst_sram_data_ok ? _GEN_10141 : _GEN_7069; // @[icache.scala 135:42]
  wire [184:0] _GEN_11166 = replace & io_inst_sram_data_ok ? _GEN_10142 : _GEN_7070; // @[icache.scala 135:42]
  wire [184:0] _GEN_11167 = replace & io_inst_sram_data_ok ? _GEN_10143 : _GEN_7071; // @[icache.scala 135:42]
  wire [184:0] _GEN_11168 = replace & io_inst_sram_data_ok ? _GEN_10144 : _GEN_7072; // @[icache.scala 135:42]
  wire [184:0] _GEN_11169 = replace & io_inst_sram_data_ok ? _GEN_10145 : _GEN_7073; // @[icache.scala 135:42]
  wire [184:0] _GEN_11170 = replace & io_inst_sram_data_ok ? _GEN_10146 : _GEN_7074; // @[icache.scala 135:42]
  wire [184:0] _GEN_11171 = replace & io_inst_sram_data_ok ? _GEN_10147 : _GEN_7075; // @[icache.scala 135:42]
  wire [184:0] _GEN_11172 = replace & io_inst_sram_data_ok ? _GEN_10148 : _GEN_7076; // @[icache.scala 135:42]
  wire [184:0] _GEN_11173 = replace & io_inst_sram_data_ok ? _GEN_10149 : _GEN_7077; // @[icache.scala 135:42]
  wire [184:0] _GEN_11174 = replace & io_inst_sram_data_ok ? _GEN_10150 : _GEN_7078; // @[icache.scala 135:42]
  wire [184:0] _GEN_11175 = replace & io_inst_sram_data_ok ? _GEN_10151 : _GEN_7079; // @[icache.scala 135:42]
  wire [184:0] _GEN_11176 = replace & io_inst_sram_data_ok ? _GEN_10152 : _GEN_7080; // @[icache.scala 135:42]
  wire [184:0] _GEN_11177 = replace & io_inst_sram_data_ok ? _GEN_10153 : _GEN_7081; // @[icache.scala 135:42]
  wire [184:0] _GEN_11178 = replace & io_inst_sram_data_ok ? _GEN_10154 : _GEN_7082; // @[icache.scala 135:42]
  wire [184:0] _GEN_11179 = replace & io_inst_sram_data_ok ? _GEN_10155 : _GEN_7083; // @[icache.scala 135:42]
  wire [184:0] _GEN_11180 = replace & io_inst_sram_data_ok ? _GEN_10156 : _GEN_7084; // @[icache.scala 135:42]
  wire [184:0] _GEN_11181 = replace & io_inst_sram_data_ok ? _GEN_10157 : _GEN_7085; // @[icache.scala 135:42]
  wire [184:0] _GEN_11182 = replace & io_inst_sram_data_ok ? _GEN_10158 : _GEN_7086; // @[icache.scala 135:42]
  wire [184:0] _GEN_11183 = replace & io_inst_sram_data_ok ? _GEN_10159 : _GEN_7087; // @[icache.scala 135:42]
  wire [184:0] _GEN_11184 = replace & io_inst_sram_data_ok ? _GEN_10160 : _GEN_7088; // @[icache.scala 135:42]
  wire [184:0] _GEN_11185 = replace & io_inst_sram_data_ok ? _GEN_10161 : _GEN_7089; // @[icache.scala 135:42]
  wire [184:0] _GEN_11186 = replace & io_inst_sram_data_ok ? _GEN_10162 : _GEN_7090; // @[icache.scala 135:42]
  wire [184:0] _GEN_11187 = replace & io_inst_sram_data_ok ? _GEN_10163 : _GEN_7091; // @[icache.scala 135:42]
  wire [184:0] _GEN_11188 = replace & io_inst_sram_data_ok ? _GEN_10164 : _GEN_7092; // @[icache.scala 135:42]
  wire [184:0] _GEN_11189 = replace & io_inst_sram_data_ok ? _GEN_10165 : _GEN_7093; // @[icache.scala 135:42]
  wire [184:0] _GEN_11190 = replace & io_inst_sram_data_ok ? _GEN_10166 : _GEN_7094; // @[icache.scala 135:42]
  wire [184:0] _GEN_11191 = replace & io_inst_sram_data_ok ? _GEN_10167 : _GEN_7095; // @[icache.scala 135:42]
  wire [184:0] _GEN_11192 = replace & io_inst_sram_data_ok ? _GEN_10168 : _GEN_7096; // @[icache.scala 135:42]
  wire [184:0] _GEN_11193 = replace & io_inst_sram_data_ok ? _GEN_10169 : _GEN_7097; // @[icache.scala 135:42]
  wire [184:0] _GEN_11194 = replace & io_inst_sram_data_ok ? _GEN_10170 : _GEN_7098; // @[icache.scala 135:42]
  wire [184:0] _GEN_11195 = replace & io_inst_sram_data_ok ? _GEN_10171 : _GEN_7099; // @[icache.scala 135:42]
  wire [184:0] _GEN_11196 = replace & io_inst_sram_data_ok ? _GEN_10172 : _GEN_7100; // @[icache.scala 135:42]
  wire [184:0] _GEN_11197 = replace & io_inst_sram_data_ok ? _GEN_10173 : _GEN_7101; // @[icache.scala 135:42]
  wire [184:0] _GEN_11198 = replace & io_inst_sram_data_ok ? _GEN_10174 : _GEN_7102; // @[icache.scala 135:42]
  wire [184:0] _GEN_11199 = replace & io_inst_sram_data_ok ? _GEN_10175 : _GEN_7103; // @[icache.scala 135:42]
  wire [184:0] _GEN_11200 = replace & io_inst_sram_data_ok ? _GEN_10176 : _GEN_7104; // @[icache.scala 135:42]
  wire [184:0] _GEN_11201 = replace & io_inst_sram_data_ok ? _GEN_10177 : _GEN_7105; // @[icache.scala 135:42]
  wire [184:0] _GEN_11202 = replace & io_inst_sram_data_ok ? _GEN_10178 : _GEN_7106; // @[icache.scala 135:42]
  wire [184:0] _GEN_11203 = replace & io_inst_sram_data_ok ? _GEN_10179 : _GEN_7107; // @[icache.scala 135:42]
  wire [184:0] _GEN_11204 = replace & io_inst_sram_data_ok ? _GEN_10180 : _GEN_7108; // @[icache.scala 135:42]
  wire [184:0] _GEN_11205 = replace & io_inst_sram_data_ok ? _GEN_10181 : _GEN_7109; // @[icache.scala 135:42]
  wire [184:0] _GEN_11206 = replace & io_inst_sram_data_ok ? _GEN_10182 : _GEN_7110; // @[icache.scala 135:42]
  wire [184:0] _GEN_11207 = replace & io_inst_sram_data_ok ? _GEN_10183 : _GEN_7111; // @[icache.scala 135:42]
  wire [184:0] _GEN_11208 = replace & io_inst_sram_data_ok ? _GEN_10184 : _GEN_7112; // @[icache.scala 135:42]
  wire [184:0] _GEN_11209 = replace & io_inst_sram_data_ok ? _GEN_10185 : _GEN_7113; // @[icache.scala 135:42]
  wire [184:0] _GEN_11210 = replace & io_inst_sram_data_ok ? _GEN_10186 : _GEN_7114; // @[icache.scala 135:42]
  wire [184:0] _GEN_11211 = replace & io_inst_sram_data_ok ? _GEN_10187 : _GEN_7115; // @[icache.scala 135:42]
  wire [184:0] _GEN_11212 = replace & io_inst_sram_data_ok ? _GEN_10188 : _GEN_7116; // @[icache.scala 135:42]
  wire [184:0] _GEN_11213 = replace & io_inst_sram_data_ok ? _GEN_10189 : _GEN_7117; // @[icache.scala 135:42]
  wire [184:0] _GEN_11214 = replace & io_inst_sram_data_ok ? _GEN_10190 : _GEN_7118; // @[icache.scala 135:42]
  wire [184:0] _GEN_11215 = replace & io_inst_sram_data_ok ? _GEN_10191 : _GEN_7119; // @[icache.scala 135:42]
  wire [184:0] _GEN_11216 = replace & io_inst_sram_data_ok ? _GEN_10192 : _GEN_7120; // @[icache.scala 135:42]
  wire [184:0] _GEN_11217 = replace & io_inst_sram_data_ok ? _GEN_10193 : _GEN_7121; // @[icache.scala 135:42]
  wire [184:0] _GEN_11218 = replace & io_inst_sram_data_ok ? _GEN_10194 : _GEN_7122; // @[icache.scala 135:42]
  wire [184:0] _GEN_11219 = replace & io_inst_sram_data_ok ? _GEN_10195 : _GEN_7123; // @[icache.scala 135:42]
  wire [184:0] _GEN_11220 = replace & io_inst_sram_data_ok ? _GEN_10196 : _GEN_7124; // @[icache.scala 135:42]
  wire [184:0] _GEN_11221 = replace & io_inst_sram_data_ok ? _GEN_10197 : _GEN_7125; // @[icache.scala 135:42]
  wire [184:0] _GEN_11222 = replace & io_inst_sram_data_ok ? _GEN_10198 : _GEN_7126; // @[icache.scala 135:42]
  wire [184:0] _GEN_11223 = replace & io_inst_sram_data_ok ? _GEN_10199 : _GEN_7127; // @[icache.scala 135:42]
  wire [184:0] _GEN_11224 = replace & io_inst_sram_data_ok ? _GEN_10200 : _GEN_7128; // @[icache.scala 135:42]
  wire [184:0] _GEN_11225 = replace & io_inst_sram_data_ok ? _GEN_10201 : _GEN_7129; // @[icache.scala 135:42]
  wire [184:0] _GEN_11226 = replace & io_inst_sram_data_ok ? _GEN_10202 : _GEN_7130; // @[icache.scala 135:42]
  wire [184:0] _GEN_11227 = replace & io_inst_sram_data_ok ? _GEN_10203 : _GEN_7131; // @[icache.scala 135:42]
  wire [184:0] _GEN_11228 = replace & io_inst_sram_data_ok ? _GEN_10204 : _GEN_7132; // @[icache.scala 135:42]
  wire [184:0] _GEN_11229 = replace & io_inst_sram_data_ok ? _GEN_10205 : _GEN_7133; // @[icache.scala 135:42]
  wire [184:0] _GEN_11230 = replace & io_inst_sram_data_ok ? _GEN_10206 : _GEN_7134; // @[icache.scala 135:42]
  wire [184:0] _GEN_11231 = replace & io_inst_sram_data_ok ? _GEN_10207 : _GEN_7135; // @[icache.scala 135:42]
  wire [184:0] _GEN_11232 = replace & io_inst_sram_data_ok ? _GEN_10208 : _GEN_7136; // @[icache.scala 135:42]
  wire [184:0] _GEN_11233 = replace & io_inst_sram_data_ok ? _GEN_10209 : _GEN_7137; // @[icache.scala 135:42]
  wire [184:0] _GEN_11234 = replace & io_inst_sram_data_ok ? _GEN_10210 : _GEN_7138; // @[icache.scala 135:42]
  wire [184:0] _GEN_11235 = replace & io_inst_sram_data_ok ? _GEN_10211 : _GEN_7139; // @[icache.scala 135:42]
  wire [184:0] _GEN_11236 = replace & io_inst_sram_data_ok ? _GEN_10212 : _GEN_7140; // @[icache.scala 135:42]
  wire [184:0] _GEN_11237 = replace & io_inst_sram_data_ok ? _GEN_10213 : _GEN_7141; // @[icache.scala 135:42]
  wire [184:0] _GEN_11238 = replace & io_inst_sram_data_ok ? _GEN_10214 : _GEN_7142; // @[icache.scala 135:42]
  wire [184:0] _GEN_11239 = replace & io_inst_sram_data_ok ? _GEN_10215 : _GEN_7143; // @[icache.scala 135:42]
  wire [184:0] _GEN_11240 = replace & io_inst_sram_data_ok ? _GEN_10216 : _GEN_7144; // @[icache.scala 135:42]
  wire [184:0] _GEN_11241 = replace & io_inst_sram_data_ok ? _GEN_10217 : _GEN_7145; // @[icache.scala 135:42]
  wire [184:0] _GEN_11242 = replace & io_inst_sram_data_ok ? _GEN_10218 : _GEN_7146; // @[icache.scala 135:42]
  wire [184:0] _GEN_11243 = replace & io_inst_sram_data_ok ? _GEN_10219 : _GEN_7147; // @[icache.scala 135:42]
  wire [184:0] _GEN_11244 = replace & io_inst_sram_data_ok ? _GEN_10220 : _GEN_7148; // @[icache.scala 135:42]
  wire [184:0] _GEN_11245 = replace & io_inst_sram_data_ok ? _GEN_10221 : _GEN_7149; // @[icache.scala 135:42]
  wire [184:0] _GEN_11246 = replace & io_inst_sram_data_ok ? _GEN_10222 : _GEN_7150; // @[icache.scala 135:42]
  wire [184:0] _GEN_11247 = replace & io_inst_sram_data_ok ? _GEN_10223 : _GEN_7151; // @[icache.scala 135:42]
  wire [184:0] _GEN_11248 = replace & io_inst_sram_data_ok ? _GEN_10224 : _GEN_7152; // @[icache.scala 135:42]
  wire [184:0] _GEN_11249 = replace & io_inst_sram_data_ok ? _GEN_10225 : _GEN_7153; // @[icache.scala 135:42]
  wire [184:0] _GEN_11250 = replace & io_inst_sram_data_ok ? _GEN_10226 : _GEN_7154; // @[icache.scala 135:42]
  wire [184:0] _GEN_11251 = replace & io_inst_sram_data_ok ? _GEN_10227 : _GEN_7155; // @[icache.scala 135:42]
  wire [184:0] _GEN_11252 = replace & io_inst_sram_data_ok ? _GEN_10228 : _GEN_7156; // @[icache.scala 135:42]
  wire [184:0] _GEN_11253 = replace & io_inst_sram_data_ok ? _GEN_10229 : _GEN_7157; // @[icache.scala 135:42]
  wire [184:0] _GEN_11254 = replace & io_inst_sram_data_ok ? _GEN_10230 : _GEN_7158; // @[icache.scala 135:42]
  wire [184:0] _GEN_11255 = replace & io_inst_sram_data_ok ? _GEN_10231 : _GEN_7159; // @[icache.scala 135:42]
  wire [184:0] _GEN_11256 = replace & io_inst_sram_data_ok ? _GEN_10232 : _GEN_7160; // @[icache.scala 135:42]
  wire [184:0] _GEN_11257 = replace & io_inst_sram_data_ok ? _GEN_10233 : _GEN_7161; // @[icache.scala 135:42]
  wire [184:0] _GEN_11258 = replace & io_inst_sram_data_ok ? _GEN_10234 : _GEN_7162; // @[icache.scala 135:42]
  wire [184:0] _GEN_11259 = replace & io_inst_sram_data_ok ? _GEN_10235 : _GEN_7163; // @[icache.scala 135:42]
  wire [184:0] _GEN_11260 = replace & io_inst_sram_data_ok ? _GEN_10236 : _GEN_7164; // @[icache.scala 135:42]
  wire [184:0] _GEN_11261 = replace & io_inst_sram_data_ok ? _GEN_10237 : _GEN_7165; // @[icache.scala 135:42]
  wire [184:0] _GEN_11262 = replace & io_inst_sram_data_ok ? _GEN_10238 : _GEN_7166; // @[icache.scala 135:42]
  wire [184:0] _GEN_11263 = replace & io_inst_sram_data_ok ? _GEN_10239 : _GEN_7167; // @[icache.scala 135:42]
  wire [184:0] _GEN_11264 = replace & io_inst_sram_data_ok ? _GEN_10240 : _GEN_7168; // @[icache.scala 135:42]
  wire [184:0] _GEN_11265 = replace & io_inst_sram_data_ok ? _GEN_10241 : _GEN_7169; // @[icache.scala 135:42]
  wire [184:0] _GEN_11266 = replace & io_inst_sram_data_ok ? _GEN_10242 : _GEN_7170; // @[icache.scala 135:42]
  wire [184:0] _GEN_11267 = replace & io_inst_sram_data_ok ? _GEN_10243 : _GEN_7171; // @[icache.scala 135:42]
  wire [184:0] _GEN_11268 = replace & io_inst_sram_data_ok ? _GEN_10244 : _GEN_7172; // @[icache.scala 135:42]
  wire [184:0] _GEN_11269 = replace & io_inst_sram_data_ok ? _GEN_10245 : _GEN_7173; // @[icache.scala 135:42]
  wire [184:0] _GEN_11270 = replace & io_inst_sram_data_ok ? _GEN_10246 : _GEN_7174; // @[icache.scala 135:42]
  wire [184:0] _GEN_11271 = replace & io_inst_sram_data_ok ? _GEN_10247 : _GEN_7175; // @[icache.scala 135:42]
  wire [184:0] _GEN_11272 = replace & io_inst_sram_data_ok ? _GEN_10248 : _GEN_7176; // @[icache.scala 135:42]
  wire [184:0] _GEN_11273 = replace & io_inst_sram_data_ok ? _GEN_10249 : _GEN_7177; // @[icache.scala 135:42]
  wire [184:0] _GEN_11274 = replace & io_inst_sram_data_ok ? _GEN_10250 : _GEN_7178; // @[icache.scala 135:42]
  wire [184:0] _GEN_11275 = replace & io_inst_sram_data_ok ? _GEN_10251 : _GEN_7179; // @[icache.scala 135:42]
  wire [184:0] _GEN_11276 = replace & io_inst_sram_data_ok ? _GEN_10252 : _GEN_7180; // @[icache.scala 135:42]
  wire [184:0] _GEN_11277 = replace & io_inst_sram_data_ok ? _GEN_10253 : _GEN_7181; // @[icache.scala 135:42]
  wire [184:0] _cache_data_T_13 = {_GEN_4095[184],1'h1,_GEN_4095[182:0]}; // @[Cat.scala 31:58]
  wire [184:0] _GEN_13326 = 10'h0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10254; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13327 = 10'h1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10255; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13328 = 10'h2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10256; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13329 = 10'h3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10257; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13330 = 10'h4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10258; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13331 = 10'h5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10259; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13332 = 10'h6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10260; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13333 = 10'h7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10261; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13334 = 10'h8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10262; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13335 = 10'h9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10263; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13336 = 10'ha == _dirty_T_1 ? _cache_data_T_13 : _GEN_10264; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13337 = 10'hb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10265; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13338 = 10'hc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10266; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13339 = 10'hd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10267; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13340 = 10'he == _dirty_T_1 ? _cache_data_T_13 : _GEN_10268; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13341 = 10'hf == _dirty_T_1 ? _cache_data_T_13 : _GEN_10269; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13342 = 10'h10 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10270; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13343 = 10'h11 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10271; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13344 = 10'h12 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10272; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13345 = 10'h13 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10273; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13346 = 10'h14 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10274; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13347 = 10'h15 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10275; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13348 = 10'h16 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10276; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13349 = 10'h17 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10277; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13350 = 10'h18 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10278; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13351 = 10'h19 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10279; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13352 = 10'h1a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10280; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13353 = 10'h1b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10281; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13354 = 10'h1c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10282; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13355 = 10'h1d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10283; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13356 = 10'h1e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10284; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13357 = 10'h1f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10285; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13358 = 10'h20 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10286; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13359 = 10'h21 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10287; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13360 = 10'h22 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10288; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13361 = 10'h23 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10289; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13362 = 10'h24 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10290; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13363 = 10'h25 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10291; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13364 = 10'h26 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10292; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13365 = 10'h27 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10293; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13366 = 10'h28 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10294; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13367 = 10'h29 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10295; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13368 = 10'h2a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10296; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13369 = 10'h2b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10297; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13370 = 10'h2c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10298; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13371 = 10'h2d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10299; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13372 = 10'h2e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10300; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13373 = 10'h2f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10301; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13374 = 10'h30 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10302; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13375 = 10'h31 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10303; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13376 = 10'h32 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10304; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13377 = 10'h33 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10305; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13378 = 10'h34 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10306; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13379 = 10'h35 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10307; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13380 = 10'h36 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10308; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13381 = 10'h37 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10309; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13382 = 10'h38 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10310; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13383 = 10'h39 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10311; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13384 = 10'h3a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10312; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13385 = 10'h3b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10313; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13386 = 10'h3c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10314; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13387 = 10'h3d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10315; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13388 = 10'h3e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10316; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13389 = 10'h3f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10317; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13390 = 10'h40 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10318; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13391 = 10'h41 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10319; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13392 = 10'h42 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10320; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13393 = 10'h43 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10321; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13394 = 10'h44 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10322; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13395 = 10'h45 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10323; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13396 = 10'h46 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10324; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13397 = 10'h47 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10325; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13398 = 10'h48 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10326; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13399 = 10'h49 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10327; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13400 = 10'h4a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10328; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13401 = 10'h4b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10329; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13402 = 10'h4c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10330; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13403 = 10'h4d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10331; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13404 = 10'h4e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10332; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13405 = 10'h4f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10333; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13406 = 10'h50 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10334; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13407 = 10'h51 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10335; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13408 = 10'h52 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10336; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13409 = 10'h53 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10337; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13410 = 10'h54 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10338; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13411 = 10'h55 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10339; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13412 = 10'h56 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10340; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13413 = 10'h57 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10341; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13414 = 10'h58 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10342; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13415 = 10'h59 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10343; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13416 = 10'h5a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10344; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13417 = 10'h5b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10345; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13418 = 10'h5c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10346; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13419 = 10'h5d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10347; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13420 = 10'h5e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10348; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13421 = 10'h5f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10349; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13422 = 10'h60 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10350; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13423 = 10'h61 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10351; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13424 = 10'h62 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10352; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13425 = 10'h63 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10353; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13426 = 10'h64 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10354; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13427 = 10'h65 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10355; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13428 = 10'h66 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10356; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13429 = 10'h67 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10357; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13430 = 10'h68 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10358; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13431 = 10'h69 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10359; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13432 = 10'h6a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10360; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13433 = 10'h6b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10361; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13434 = 10'h6c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10362; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13435 = 10'h6d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10363; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13436 = 10'h6e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10364; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13437 = 10'h6f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10365; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13438 = 10'h70 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10366; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13439 = 10'h71 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10367; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13440 = 10'h72 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10368; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13441 = 10'h73 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10369; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13442 = 10'h74 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10370; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13443 = 10'h75 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10371; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13444 = 10'h76 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10372; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13445 = 10'h77 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10373; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13446 = 10'h78 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10374; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13447 = 10'h79 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10375; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13448 = 10'h7a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10376; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13449 = 10'h7b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10377; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13450 = 10'h7c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10378; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13451 = 10'h7d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10379; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13452 = 10'h7e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10380; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13453 = 10'h7f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10381; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13454 = 10'h80 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10382; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13455 = 10'h81 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10383; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13456 = 10'h82 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10384; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13457 = 10'h83 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10385; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13458 = 10'h84 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10386; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13459 = 10'h85 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10387; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13460 = 10'h86 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10388; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13461 = 10'h87 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10389; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13462 = 10'h88 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10390; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13463 = 10'h89 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10391; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13464 = 10'h8a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10392; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13465 = 10'h8b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10393; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13466 = 10'h8c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10394; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13467 = 10'h8d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10395; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13468 = 10'h8e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10396; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13469 = 10'h8f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10397; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13470 = 10'h90 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10398; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13471 = 10'h91 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10399; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13472 = 10'h92 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10400; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13473 = 10'h93 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10401; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13474 = 10'h94 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10402; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13475 = 10'h95 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10403; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13476 = 10'h96 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10404; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13477 = 10'h97 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10405; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13478 = 10'h98 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10406; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13479 = 10'h99 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10407; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13480 = 10'h9a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10408; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13481 = 10'h9b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10409; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13482 = 10'h9c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10410; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13483 = 10'h9d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10411; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13484 = 10'h9e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10412; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13485 = 10'h9f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10413; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13486 = 10'ha0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10414; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13487 = 10'ha1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10415; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13488 = 10'ha2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10416; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13489 = 10'ha3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10417; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13490 = 10'ha4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10418; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13491 = 10'ha5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10419; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13492 = 10'ha6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10420; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13493 = 10'ha7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10421; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13494 = 10'ha8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10422; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13495 = 10'ha9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10423; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13496 = 10'haa == _dirty_T_1 ? _cache_data_T_13 : _GEN_10424; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13497 = 10'hab == _dirty_T_1 ? _cache_data_T_13 : _GEN_10425; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13498 = 10'hac == _dirty_T_1 ? _cache_data_T_13 : _GEN_10426; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13499 = 10'had == _dirty_T_1 ? _cache_data_T_13 : _GEN_10427; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13500 = 10'hae == _dirty_T_1 ? _cache_data_T_13 : _GEN_10428; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13501 = 10'haf == _dirty_T_1 ? _cache_data_T_13 : _GEN_10429; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13502 = 10'hb0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10430; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13503 = 10'hb1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10431; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13504 = 10'hb2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10432; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13505 = 10'hb3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10433; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13506 = 10'hb4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10434; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13507 = 10'hb5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10435; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13508 = 10'hb6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10436; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13509 = 10'hb7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10437; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13510 = 10'hb8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10438; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13511 = 10'hb9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10439; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13512 = 10'hba == _dirty_T_1 ? _cache_data_T_13 : _GEN_10440; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13513 = 10'hbb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10441; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13514 = 10'hbc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10442; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13515 = 10'hbd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10443; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13516 = 10'hbe == _dirty_T_1 ? _cache_data_T_13 : _GEN_10444; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13517 = 10'hbf == _dirty_T_1 ? _cache_data_T_13 : _GEN_10445; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13518 = 10'hc0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10446; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13519 = 10'hc1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10447; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13520 = 10'hc2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10448; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13521 = 10'hc3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10449; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13522 = 10'hc4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10450; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13523 = 10'hc5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10451; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13524 = 10'hc6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10452; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13525 = 10'hc7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10453; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13526 = 10'hc8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10454; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13527 = 10'hc9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10455; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13528 = 10'hca == _dirty_T_1 ? _cache_data_T_13 : _GEN_10456; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13529 = 10'hcb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10457; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13530 = 10'hcc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10458; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13531 = 10'hcd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10459; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13532 = 10'hce == _dirty_T_1 ? _cache_data_T_13 : _GEN_10460; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13533 = 10'hcf == _dirty_T_1 ? _cache_data_T_13 : _GEN_10461; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13534 = 10'hd0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10462; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13535 = 10'hd1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10463; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13536 = 10'hd2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10464; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13537 = 10'hd3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10465; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13538 = 10'hd4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10466; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13539 = 10'hd5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10467; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13540 = 10'hd6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10468; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13541 = 10'hd7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10469; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13542 = 10'hd8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10470; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13543 = 10'hd9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10471; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13544 = 10'hda == _dirty_T_1 ? _cache_data_T_13 : _GEN_10472; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13545 = 10'hdb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10473; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13546 = 10'hdc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10474; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13547 = 10'hdd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10475; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13548 = 10'hde == _dirty_T_1 ? _cache_data_T_13 : _GEN_10476; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13549 = 10'hdf == _dirty_T_1 ? _cache_data_T_13 : _GEN_10477; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13550 = 10'he0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10478; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13551 = 10'he1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10479; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13552 = 10'he2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10480; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13553 = 10'he3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10481; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13554 = 10'he4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10482; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13555 = 10'he5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10483; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13556 = 10'he6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10484; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13557 = 10'he7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10485; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13558 = 10'he8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10486; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13559 = 10'he9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10487; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13560 = 10'hea == _dirty_T_1 ? _cache_data_T_13 : _GEN_10488; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13561 = 10'heb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10489; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13562 = 10'hec == _dirty_T_1 ? _cache_data_T_13 : _GEN_10490; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13563 = 10'hed == _dirty_T_1 ? _cache_data_T_13 : _GEN_10491; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13564 = 10'hee == _dirty_T_1 ? _cache_data_T_13 : _GEN_10492; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13565 = 10'hef == _dirty_T_1 ? _cache_data_T_13 : _GEN_10493; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13566 = 10'hf0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10494; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13567 = 10'hf1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10495; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13568 = 10'hf2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10496; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13569 = 10'hf3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10497; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13570 = 10'hf4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10498; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13571 = 10'hf5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10499; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13572 = 10'hf6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10500; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13573 = 10'hf7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10501; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13574 = 10'hf8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10502; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13575 = 10'hf9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10503; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13576 = 10'hfa == _dirty_T_1 ? _cache_data_T_13 : _GEN_10504; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13577 = 10'hfb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10505; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13578 = 10'hfc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10506; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13579 = 10'hfd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10507; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13580 = 10'hfe == _dirty_T_1 ? _cache_data_T_13 : _GEN_10508; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13581 = 10'hff == _dirty_T_1 ? _cache_data_T_13 : _GEN_10509; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13582 = 10'h100 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10510; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13583 = 10'h101 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10511; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13584 = 10'h102 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10512; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13585 = 10'h103 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10513; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13586 = 10'h104 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10514; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13587 = 10'h105 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10515; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13588 = 10'h106 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10516; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13589 = 10'h107 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10517; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13590 = 10'h108 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10518; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13591 = 10'h109 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10519; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13592 = 10'h10a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10520; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13593 = 10'h10b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10521; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13594 = 10'h10c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10522; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13595 = 10'h10d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10523; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13596 = 10'h10e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10524; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13597 = 10'h10f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10525; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13598 = 10'h110 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10526; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13599 = 10'h111 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10527; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13600 = 10'h112 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10528; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13601 = 10'h113 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10529; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13602 = 10'h114 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10530; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13603 = 10'h115 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10531; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13604 = 10'h116 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10532; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13605 = 10'h117 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10533; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13606 = 10'h118 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10534; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13607 = 10'h119 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10535; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13608 = 10'h11a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10536; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13609 = 10'h11b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10537; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13610 = 10'h11c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10538; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13611 = 10'h11d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10539; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13612 = 10'h11e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10540; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13613 = 10'h11f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10541; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13614 = 10'h120 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10542; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13615 = 10'h121 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10543; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13616 = 10'h122 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10544; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13617 = 10'h123 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10545; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13618 = 10'h124 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10546; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13619 = 10'h125 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10547; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13620 = 10'h126 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10548; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13621 = 10'h127 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10549; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13622 = 10'h128 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10550; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13623 = 10'h129 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10551; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13624 = 10'h12a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10552; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13625 = 10'h12b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10553; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13626 = 10'h12c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10554; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13627 = 10'h12d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10555; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13628 = 10'h12e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10556; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13629 = 10'h12f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10557; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13630 = 10'h130 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10558; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13631 = 10'h131 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10559; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13632 = 10'h132 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10560; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13633 = 10'h133 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10561; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13634 = 10'h134 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10562; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13635 = 10'h135 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10563; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13636 = 10'h136 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10564; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13637 = 10'h137 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10565; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13638 = 10'h138 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10566; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13639 = 10'h139 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10567; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13640 = 10'h13a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10568; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13641 = 10'h13b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10569; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13642 = 10'h13c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10570; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13643 = 10'h13d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10571; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13644 = 10'h13e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10572; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13645 = 10'h13f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10573; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13646 = 10'h140 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10574; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13647 = 10'h141 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10575; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13648 = 10'h142 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10576; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13649 = 10'h143 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10577; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13650 = 10'h144 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10578; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13651 = 10'h145 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10579; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13652 = 10'h146 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10580; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13653 = 10'h147 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10581; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13654 = 10'h148 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10582; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13655 = 10'h149 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10583; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13656 = 10'h14a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10584; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13657 = 10'h14b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10585; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13658 = 10'h14c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10586; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13659 = 10'h14d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10587; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13660 = 10'h14e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10588; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13661 = 10'h14f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10589; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13662 = 10'h150 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10590; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13663 = 10'h151 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10591; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13664 = 10'h152 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10592; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13665 = 10'h153 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10593; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13666 = 10'h154 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10594; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13667 = 10'h155 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10595; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13668 = 10'h156 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10596; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13669 = 10'h157 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10597; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13670 = 10'h158 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10598; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13671 = 10'h159 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10599; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13672 = 10'h15a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10600; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13673 = 10'h15b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10601; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13674 = 10'h15c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10602; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13675 = 10'h15d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10603; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13676 = 10'h15e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10604; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13677 = 10'h15f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10605; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13678 = 10'h160 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10606; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13679 = 10'h161 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10607; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13680 = 10'h162 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10608; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13681 = 10'h163 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10609; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13682 = 10'h164 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10610; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13683 = 10'h165 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10611; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13684 = 10'h166 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10612; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13685 = 10'h167 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10613; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13686 = 10'h168 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10614; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13687 = 10'h169 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10615; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13688 = 10'h16a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10616; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13689 = 10'h16b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10617; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13690 = 10'h16c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10618; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13691 = 10'h16d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10619; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13692 = 10'h16e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10620; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13693 = 10'h16f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10621; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13694 = 10'h170 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10622; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13695 = 10'h171 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10623; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13696 = 10'h172 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10624; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13697 = 10'h173 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10625; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13698 = 10'h174 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10626; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13699 = 10'h175 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10627; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13700 = 10'h176 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10628; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13701 = 10'h177 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10629; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13702 = 10'h178 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10630; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13703 = 10'h179 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10631; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13704 = 10'h17a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10632; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13705 = 10'h17b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10633; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13706 = 10'h17c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10634; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13707 = 10'h17d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10635; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13708 = 10'h17e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10636; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13709 = 10'h17f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10637; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13710 = 10'h180 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10638; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13711 = 10'h181 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10639; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13712 = 10'h182 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10640; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13713 = 10'h183 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10641; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13714 = 10'h184 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10642; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13715 = 10'h185 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10643; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13716 = 10'h186 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10644; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13717 = 10'h187 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10645; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13718 = 10'h188 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10646; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13719 = 10'h189 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10647; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13720 = 10'h18a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10648; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13721 = 10'h18b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10649; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13722 = 10'h18c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10650; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13723 = 10'h18d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10651; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13724 = 10'h18e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10652; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13725 = 10'h18f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10653; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13726 = 10'h190 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10654; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13727 = 10'h191 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10655; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13728 = 10'h192 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10656; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13729 = 10'h193 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10657; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13730 = 10'h194 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10658; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13731 = 10'h195 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10659; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13732 = 10'h196 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10660; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13733 = 10'h197 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10661; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13734 = 10'h198 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10662; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13735 = 10'h199 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10663; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13736 = 10'h19a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10664; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13737 = 10'h19b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10665; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13738 = 10'h19c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10666; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13739 = 10'h19d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10667; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13740 = 10'h19e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10668; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13741 = 10'h19f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10669; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13742 = 10'h1a0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10670; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13743 = 10'h1a1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10671; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13744 = 10'h1a2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10672; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13745 = 10'h1a3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10673; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13746 = 10'h1a4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10674; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13747 = 10'h1a5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10675; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13748 = 10'h1a6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10676; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13749 = 10'h1a7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10677; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13750 = 10'h1a8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10678; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13751 = 10'h1a9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10679; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13752 = 10'h1aa == _dirty_T_1 ? _cache_data_T_13 : _GEN_10680; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13753 = 10'h1ab == _dirty_T_1 ? _cache_data_T_13 : _GEN_10681; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13754 = 10'h1ac == _dirty_T_1 ? _cache_data_T_13 : _GEN_10682; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13755 = 10'h1ad == _dirty_T_1 ? _cache_data_T_13 : _GEN_10683; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13756 = 10'h1ae == _dirty_T_1 ? _cache_data_T_13 : _GEN_10684; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13757 = 10'h1af == _dirty_T_1 ? _cache_data_T_13 : _GEN_10685; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13758 = 10'h1b0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10686; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13759 = 10'h1b1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10687; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13760 = 10'h1b2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10688; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13761 = 10'h1b3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10689; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13762 = 10'h1b4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10690; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13763 = 10'h1b5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10691; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13764 = 10'h1b6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10692; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13765 = 10'h1b7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10693; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13766 = 10'h1b8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10694; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13767 = 10'h1b9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10695; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13768 = 10'h1ba == _dirty_T_1 ? _cache_data_T_13 : _GEN_10696; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13769 = 10'h1bb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10697; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13770 = 10'h1bc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10698; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13771 = 10'h1bd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10699; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13772 = 10'h1be == _dirty_T_1 ? _cache_data_T_13 : _GEN_10700; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13773 = 10'h1bf == _dirty_T_1 ? _cache_data_T_13 : _GEN_10701; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13774 = 10'h1c0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10702; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13775 = 10'h1c1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10703; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13776 = 10'h1c2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10704; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13777 = 10'h1c3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10705; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13778 = 10'h1c4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10706; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13779 = 10'h1c5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10707; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13780 = 10'h1c6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10708; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13781 = 10'h1c7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10709; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13782 = 10'h1c8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10710; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13783 = 10'h1c9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10711; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13784 = 10'h1ca == _dirty_T_1 ? _cache_data_T_13 : _GEN_10712; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13785 = 10'h1cb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10713; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13786 = 10'h1cc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10714; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13787 = 10'h1cd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10715; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13788 = 10'h1ce == _dirty_T_1 ? _cache_data_T_13 : _GEN_10716; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13789 = 10'h1cf == _dirty_T_1 ? _cache_data_T_13 : _GEN_10717; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13790 = 10'h1d0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10718; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13791 = 10'h1d1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10719; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13792 = 10'h1d2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10720; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13793 = 10'h1d3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10721; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13794 = 10'h1d4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10722; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13795 = 10'h1d5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10723; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13796 = 10'h1d6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10724; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13797 = 10'h1d7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10725; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13798 = 10'h1d8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10726; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13799 = 10'h1d9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10727; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13800 = 10'h1da == _dirty_T_1 ? _cache_data_T_13 : _GEN_10728; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13801 = 10'h1db == _dirty_T_1 ? _cache_data_T_13 : _GEN_10729; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13802 = 10'h1dc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10730; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13803 = 10'h1dd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10731; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13804 = 10'h1de == _dirty_T_1 ? _cache_data_T_13 : _GEN_10732; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13805 = 10'h1df == _dirty_T_1 ? _cache_data_T_13 : _GEN_10733; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13806 = 10'h1e0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10734; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13807 = 10'h1e1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10735; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13808 = 10'h1e2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10736; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13809 = 10'h1e3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10737; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13810 = 10'h1e4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10738; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13811 = 10'h1e5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10739; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13812 = 10'h1e6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10740; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13813 = 10'h1e7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10741; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13814 = 10'h1e8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10742; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13815 = 10'h1e9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10743; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13816 = 10'h1ea == _dirty_T_1 ? _cache_data_T_13 : _GEN_10744; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13817 = 10'h1eb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10745; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13818 = 10'h1ec == _dirty_T_1 ? _cache_data_T_13 : _GEN_10746; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13819 = 10'h1ed == _dirty_T_1 ? _cache_data_T_13 : _GEN_10747; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13820 = 10'h1ee == _dirty_T_1 ? _cache_data_T_13 : _GEN_10748; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13821 = 10'h1ef == _dirty_T_1 ? _cache_data_T_13 : _GEN_10749; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13822 = 10'h1f0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10750; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13823 = 10'h1f1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10751; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13824 = 10'h1f2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10752; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13825 = 10'h1f3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10753; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13826 = 10'h1f4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10754; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13827 = 10'h1f5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10755; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13828 = 10'h1f6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10756; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13829 = 10'h1f7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10757; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13830 = 10'h1f8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10758; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13831 = 10'h1f9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10759; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13832 = 10'h1fa == _dirty_T_1 ? _cache_data_T_13 : _GEN_10760; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13833 = 10'h1fb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10761; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13834 = 10'h1fc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10762; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13835 = 10'h1fd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10763; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13836 = 10'h1fe == _dirty_T_1 ? _cache_data_T_13 : _GEN_10764; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13837 = 10'h1ff == _dirty_T_1 ? _cache_data_T_13 : _GEN_10765; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13838 = 10'h200 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10766; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13839 = 10'h201 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10767; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13840 = 10'h202 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10768; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13841 = 10'h203 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10769; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13842 = 10'h204 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10770; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13843 = 10'h205 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10771; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13844 = 10'h206 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10772; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13845 = 10'h207 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10773; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13846 = 10'h208 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10774; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13847 = 10'h209 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10775; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13848 = 10'h20a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10776; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13849 = 10'h20b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10777; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13850 = 10'h20c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10778; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13851 = 10'h20d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10779; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13852 = 10'h20e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10780; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13853 = 10'h20f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10781; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13854 = 10'h210 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10782; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13855 = 10'h211 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10783; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13856 = 10'h212 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10784; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13857 = 10'h213 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10785; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13858 = 10'h214 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10786; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13859 = 10'h215 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10787; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13860 = 10'h216 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10788; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13861 = 10'h217 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10789; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13862 = 10'h218 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10790; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13863 = 10'h219 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10791; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13864 = 10'h21a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10792; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13865 = 10'h21b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10793; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13866 = 10'h21c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10794; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13867 = 10'h21d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10795; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13868 = 10'h21e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10796; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13869 = 10'h21f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10797; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13870 = 10'h220 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10798; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13871 = 10'h221 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10799; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13872 = 10'h222 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10800; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13873 = 10'h223 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10801; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13874 = 10'h224 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10802; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13875 = 10'h225 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10803; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13876 = 10'h226 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10804; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13877 = 10'h227 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10805; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13878 = 10'h228 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10806; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13879 = 10'h229 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10807; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13880 = 10'h22a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10808; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13881 = 10'h22b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10809; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13882 = 10'h22c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10810; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13883 = 10'h22d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10811; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13884 = 10'h22e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10812; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13885 = 10'h22f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10813; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13886 = 10'h230 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10814; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13887 = 10'h231 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10815; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13888 = 10'h232 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10816; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13889 = 10'h233 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10817; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13890 = 10'h234 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10818; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13891 = 10'h235 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10819; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13892 = 10'h236 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10820; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13893 = 10'h237 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10821; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13894 = 10'h238 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10822; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13895 = 10'h239 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10823; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13896 = 10'h23a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10824; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13897 = 10'h23b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10825; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13898 = 10'h23c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10826; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13899 = 10'h23d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10827; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13900 = 10'h23e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10828; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13901 = 10'h23f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10829; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13902 = 10'h240 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10830; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13903 = 10'h241 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10831; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13904 = 10'h242 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10832; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13905 = 10'h243 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10833; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13906 = 10'h244 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10834; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13907 = 10'h245 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10835; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13908 = 10'h246 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10836; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13909 = 10'h247 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10837; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13910 = 10'h248 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10838; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13911 = 10'h249 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10839; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13912 = 10'h24a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10840; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13913 = 10'h24b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10841; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13914 = 10'h24c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10842; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13915 = 10'h24d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10843; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13916 = 10'h24e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10844; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13917 = 10'h24f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10845; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13918 = 10'h250 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10846; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13919 = 10'h251 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10847; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13920 = 10'h252 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10848; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13921 = 10'h253 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10849; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13922 = 10'h254 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10850; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13923 = 10'h255 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10851; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13924 = 10'h256 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10852; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13925 = 10'h257 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10853; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13926 = 10'h258 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10854; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13927 = 10'h259 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10855; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13928 = 10'h25a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10856; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13929 = 10'h25b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10857; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13930 = 10'h25c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10858; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13931 = 10'h25d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10859; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13932 = 10'h25e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10860; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13933 = 10'h25f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10861; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13934 = 10'h260 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10862; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13935 = 10'h261 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10863; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13936 = 10'h262 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10864; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13937 = 10'h263 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10865; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13938 = 10'h264 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10866; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13939 = 10'h265 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10867; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13940 = 10'h266 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10868; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13941 = 10'h267 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10869; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13942 = 10'h268 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10870; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13943 = 10'h269 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10871; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13944 = 10'h26a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10872; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13945 = 10'h26b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10873; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13946 = 10'h26c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10874; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13947 = 10'h26d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10875; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13948 = 10'h26e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10876; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13949 = 10'h26f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10877; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13950 = 10'h270 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10878; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13951 = 10'h271 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10879; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13952 = 10'h272 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10880; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13953 = 10'h273 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10881; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13954 = 10'h274 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10882; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13955 = 10'h275 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10883; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13956 = 10'h276 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10884; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13957 = 10'h277 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10885; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13958 = 10'h278 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10886; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13959 = 10'h279 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10887; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13960 = 10'h27a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10888; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13961 = 10'h27b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10889; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13962 = 10'h27c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10890; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13963 = 10'h27d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10891; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13964 = 10'h27e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10892; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13965 = 10'h27f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10893; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13966 = 10'h280 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10894; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13967 = 10'h281 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10895; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13968 = 10'h282 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10896; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13969 = 10'h283 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10897; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13970 = 10'h284 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10898; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13971 = 10'h285 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10899; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13972 = 10'h286 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10900; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13973 = 10'h287 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10901; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13974 = 10'h288 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10902; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13975 = 10'h289 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10903; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13976 = 10'h28a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10904; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13977 = 10'h28b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10905; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13978 = 10'h28c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10906; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13979 = 10'h28d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10907; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13980 = 10'h28e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10908; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13981 = 10'h28f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10909; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13982 = 10'h290 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10910; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13983 = 10'h291 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10911; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13984 = 10'h292 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10912; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13985 = 10'h293 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10913; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13986 = 10'h294 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10914; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13987 = 10'h295 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10915; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13988 = 10'h296 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10916; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13989 = 10'h297 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10917; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13990 = 10'h298 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10918; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13991 = 10'h299 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10919; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13992 = 10'h29a == _dirty_T_1 ? _cache_data_T_13 : _GEN_10920; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13993 = 10'h29b == _dirty_T_1 ? _cache_data_T_13 : _GEN_10921; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13994 = 10'h29c == _dirty_T_1 ? _cache_data_T_13 : _GEN_10922; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13995 = 10'h29d == _dirty_T_1 ? _cache_data_T_13 : _GEN_10923; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13996 = 10'h29e == _dirty_T_1 ? _cache_data_T_13 : _GEN_10924; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13997 = 10'h29f == _dirty_T_1 ? _cache_data_T_13 : _GEN_10925; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13998 = 10'h2a0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10926; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_13999 = 10'h2a1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10927; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14000 = 10'h2a2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10928; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14001 = 10'h2a3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10929; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14002 = 10'h2a4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10930; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14003 = 10'h2a5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10931; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14004 = 10'h2a6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10932; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14005 = 10'h2a7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10933; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14006 = 10'h2a8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10934; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14007 = 10'h2a9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10935; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14008 = 10'h2aa == _dirty_T_1 ? _cache_data_T_13 : _GEN_10936; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14009 = 10'h2ab == _dirty_T_1 ? _cache_data_T_13 : _GEN_10937; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14010 = 10'h2ac == _dirty_T_1 ? _cache_data_T_13 : _GEN_10938; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14011 = 10'h2ad == _dirty_T_1 ? _cache_data_T_13 : _GEN_10939; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14012 = 10'h2ae == _dirty_T_1 ? _cache_data_T_13 : _GEN_10940; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14013 = 10'h2af == _dirty_T_1 ? _cache_data_T_13 : _GEN_10941; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14014 = 10'h2b0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10942; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14015 = 10'h2b1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10943; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14016 = 10'h2b2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10944; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14017 = 10'h2b3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10945; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14018 = 10'h2b4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10946; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14019 = 10'h2b5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10947; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14020 = 10'h2b6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10948; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14021 = 10'h2b7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10949; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14022 = 10'h2b8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10950; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14023 = 10'h2b9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10951; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14024 = 10'h2ba == _dirty_T_1 ? _cache_data_T_13 : _GEN_10952; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14025 = 10'h2bb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10953; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14026 = 10'h2bc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10954; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14027 = 10'h2bd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10955; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14028 = 10'h2be == _dirty_T_1 ? _cache_data_T_13 : _GEN_10956; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14029 = 10'h2bf == _dirty_T_1 ? _cache_data_T_13 : _GEN_10957; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14030 = 10'h2c0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10958; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14031 = 10'h2c1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10959; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14032 = 10'h2c2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10960; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14033 = 10'h2c3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10961; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14034 = 10'h2c4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10962; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14035 = 10'h2c5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10963; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14036 = 10'h2c6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10964; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14037 = 10'h2c7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10965; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14038 = 10'h2c8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10966; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14039 = 10'h2c9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10967; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14040 = 10'h2ca == _dirty_T_1 ? _cache_data_T_13 : _GEN_10968; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14041 = 10'h2cb == _dirty_T_1 ? _cache_data_T_13 : _GEN_10969; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14042 = 10'h2cc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10970; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14043 = 10'h2cd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10971; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14044 = 10'h2ce == _dirty_T_1 ? _cache_data_T_13 : _GEN_10972; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14045 = 10'h2cf == _dirty_T_1 ? _cache_data_T_13 : _GEN_10973; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14046 = 10'h2d0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10974; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14047 = 10'h2d1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10975; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14048 = 10'h2d2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10976; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14049 = 10'h2d3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10977; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14050 = 10'h2d4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10978; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14051 = 10'h2d5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10979; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14052 = 10'h2d6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10980; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14053 = 10'h2d7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10981; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14054 = 10'h2d8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10982; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14055 = 10'h2d9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10983; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14056 = 10'h2da == _dirty_T_1 ? _cache_data_T_13 : _GEN_10984; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14057 = 10'h2db == _dirty_T_1 ? _cache_data_T_13 : _GEN_10985; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14058 = 10'h2dc == _dirty_T_1 ? _cache_data_T_13 : _GEN_10986; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14059 = 10'h2dd == _dirty_T_1 ? _cache_data_T_13 : _GEN_10987; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14060 = 10'h2de == _dirty_T_1 ? _cache_data_T_13 : _GEN_10988; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14061 = 10'h2df == _dirty_T_1 ? _cache_data_T_13 : _GEN_10989; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14062 = 10'h2e0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10990; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14063 = 10'h2e1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10991; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14064 = 10'h2e2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10992; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14065 = 10'h2e3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10993; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14066 = 10'h2e4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10994; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14067 = 10'h2e5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10995; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14068 = 10'h2e6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10996; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14069 = 10'h2e7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10997; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14070 = 10'h2e8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10998; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14071 = 10'h2e9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_10999; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14072 = 10'h2ea == _dirty_T_1 ? _cache_data_T_13 : _GEN_11000; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14073 = 10'h2eb == _dirty_T_1 ? _cache_data_T_13 : _GEN_11001; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14074 = 10'h2ec == _dirty_T_1 ? _cache_data_T_13 : _GEN_11002; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14075 = 10'h2ed == _dirty_T_1 ? _cache_data_T_13 : _GEN_11003; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14076 = 10'h2ee == _dirty_T_1 ? _cache_data_T_13 : _GEN_11004; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14077 = 10'h2ef == _dirty_T_1 ? _cache_data_T_13 : _GEN_11005; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14078 = 10'h2f0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11006; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14079 = 10'h2f1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11007; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14080 = 10'h2f2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11008; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14081 = 10'h2f3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11009; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14082 = 10'h2f4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11010; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14083 = 10'h2f5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11011; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14084 = 10'h2f6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11012; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14085 = 10'h2f7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11013; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14086 = 10'h2f8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11014; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14087 = 10'h2f9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11015; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14088 = 10'h2fa == _dirty_T_1 ? _cache_data_T_13 : _GEN_11016; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14089 = 10'h2fb == _dirty_T_1 ? _cache_data_T_13 : _GEN_11017; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14090 = 10'h2fc == _dirty_T_1 ? _cache_data_T_13 : _GEN_11018; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14091 = 10'h2fd == _dirty_T_1 ? _cache_data_T_13 : _GEN_11019; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14092 = 10'h2fe == _dirty_T_1 ? _cache_data_T_13 : _GEN_11020; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14093 = 10'h2ff == _dirty_T_1 ? _cache_data_T_13 : _GEN_11021; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14094 = 10'h300 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11022; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14095 = 10'h301 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11023; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14096 = 10'h302 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11024; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14097 = 10'h303 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11025; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14098 = 10'h304 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11026; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14099 = 10'h305 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11027; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14100 = 10'h306 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11028; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14101 = 10'h307 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11029; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14102 = 10'h308 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11030; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14103 = 10'h309 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11031; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14104 = 10'h30a == _dirty_T_1 ? _cache_data_T_13 : _GEN_11032; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14105 = 10'h30b == _dirty_T_1 ? _cache_data_T_13 : _GEN_11033; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14106 = 10'h30c == _dirty_T_1 ? _cache_data_T_13 : _GEN_11034; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14107 = 10'h30d == _dirty_T_1 ? _cache_data_T_13 : _GEN_11035; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14108 = 10'h30e == _dirty_T_1 ? _cache_data_T_13 : _GEN_11036; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14109 = 10'h30f == _dirty_T_1 ? _cache_data_T_13 : _GEN_11037; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14110 = 10'h310 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11038; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14111 = 10'h311 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11039; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14112 = 10'h312 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11040; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14113 = 10'h313 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11041; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14114 = 10'h314 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11042; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14115 = 10'h315 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11043; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14116 = 10'h316 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11044; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14117 = 10'h317 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11045; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14118 = 10'h318 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11046; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14119 = 10'h319 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11047; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14120 = 10'h31a == _dirty_T_1 ? _cache_data_T_13 : _GEN_11048; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14121 = 10'h31b == _dirty_T_1 ? _cache_data_T_13 : _GEN_11049; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14122 = 10'h31c == _dirty_T_1 ? _cache_data_T_13 : _GEN_11050; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14123 = 10'h31d == _dirty_T_1 ? _cache_data_T_13 : _GEN_11051; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14124 = 10'h31e == _dirty_T_1 ? _cache_data_T_13 : _GEN_11052; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14125 = 10'h31f == _dirty_T_1 ? _cache_data_T_13 : _GEN_11053; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14126 = 10'h320 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11054; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14127 = 10'h321 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11055; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14128 = 10'h322 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11056; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14129 = 10'h323 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11057; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14130 = 10'h324 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11058; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14131 = 10'h325 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11059; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14132 = 10'h326 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11060; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14133 = 10'h327 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11061; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14134 = 10'h328 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11062; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14135 = 10'h329 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11063; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14136 = 10'h32a == _dirty_T_1 ? _cache_data_T_13 : _GEN_11064; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14137 = 10'h32b == _dirty_T_1 ? _cache_data_T_13 : _GEN_11065; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14138 = 10'h32c == _dirty_T_1 ? _cache_data_T_13 : _GEN_11066; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14139 = 10'h32d == _dirty_T_1 ? _cache_data_T_13 : _GEN_11067; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14140 = 10'h32e == _dirty_T_1 ? _cache_data_T_13 : _GEN_11068; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14141 = 10'h32f == _dirty_T_1 ? _cache_data_T_13 : _GEN_11069; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14142 = 10'h330 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11070; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14143 = 10'h331 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11071; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14144 = 10'h332 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11072; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14145 = 10'h333 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11073; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14146 = 10'h334 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11074; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14147 = 10'h335 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11075; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14148 = 10'h336 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11076; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14149 = 10'h337 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11077; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14150 = 10'h338 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11078; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14151 = 10'h339 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11079; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14152 = 10'h33a == _dirty_T_1 ? _cache_data_T_13 : _GEN_11080; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14153 = 10'h33b == _dirty_T_1 ? _cache_data_T_13 : _GEN_11081; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14154 = 10'h33c == _dirty_T_1 ? _cache_data_T_13 : _GEN_11082; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14155 = 10'h33d == _dirty_T_1 ? _cache_data_T_13 : _GEN_11083; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14156 = 10'h33e == _dirty_T_1 ? _cache_data_T_13 : _GEN_11084; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14157 = 10'h33f == _dirty_T_1 ? _cache_data_T_13 : _GEN_11085; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14158 = 10'h340 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11086; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14159 = 10'h341 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11087; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14160 = 10'h342 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11088; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14161 = 10'h343 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11089; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14162 = 10'h344 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11090; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14163 = 10'h345 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11091; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14164 = 10'h346 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11092; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14165 = 10'h347 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11093; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14166 = 10'h348 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11094; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14167 = 10'h349 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11095; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14168 = 10'h34a == _dirty_T_1 ? _cache_data_T_13 : _GEN_11096; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14169 = 10'h34b == _dirty_T_1 ? _cache_data_T_13 : _GEN_11097; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14170 = 10'h34c == _dirty_T_1 ? _cache_data_T_13 : _GEN_11098; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14171 = 10'h34d == _dirty_T_1 ? _cache_data_T_13 : _GEN_11099; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14172 = 10'h34e == _dirty_T_1 ? _cache_data_T_13 : _GEN_11100; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14173 = 10'h34f == _dirty_T_1 ? _cache_data_T_13 : _GEN_11101; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14174 = 10'h350 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11102; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14175 = 10'h351 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11103; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14176 = 10'h352 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11104; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14177 = 10'h353 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11105; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14178 = 10'h354 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11106; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14179 = 10'h355 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11107; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14180 = 10'h356 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11108; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14181 = 10'h357 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11109; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14182 = 10'h358 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11110; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14183 = 10'h359 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11111; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14184 = 10'h35a == _dirty_T_1 ? _cache_data_T_13 : _GEN_11112; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14185 = 10'h35b == _dirty_T_1 ? _cache_data_T_13 : _GEN_11113; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14186 = 10'h35c == _dirty_T_1 ? _cache_data_T_13 : _GEN_11114; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14187 = 10'h35d == _dirty_T_1 ? _cache_data_T_13 : _GEN_11115; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14188 = 10'h35e == _dirty_T_1 ? _cache_data_T_13 : _GEN_11116; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14189 = 10'h35f == _dirty_T_1 ? _cache_data_T_13 : _GEN_11117; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14190 = 10'h360 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11118; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14191 = 10'h361 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11119; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14192 = 10'h362 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11120; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14193 = 10'h363 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11121; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14194 = 10'h364 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11122; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14195 = 10'h365 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11123; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14196 = 10'h366 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11124; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14197 = 10'h367 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11125; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14198 = 10'h368 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11126; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14199 = 10'h369 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11127; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14200 = 10'h36a == _dirty_T_1 ? _cache_data_T_13 : _GEN_11128; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14201 = 10'h36b == _dirty_T_1 ? _cache_data_T_13 : _GEN_11129; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14202 = 10'h36c == _dirty_T_1 ? _cache_data_T_13 : _GEN_11130; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14203 = 10'h36d == _dirty_T_1 ? _cache_data_T_13 : _GEN_11131; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14204 = 10'h36e == _dirty_T_1 ? _cache_data_T_13 : _GEN_11132; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14205 = 10'h36f == _dirty_T_1 ? _cache_data_T_13 : _GEN_11133; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14206 = 10'h370 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11134; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14207 = 10'h371 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11135; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14208 = 10'h372 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11136; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14209 = 10'h373 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11137; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14210 = 10'h374 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11138; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14211 = 10'h375 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11139; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14212 = 10'h376 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11140; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14213 = 10'h377 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11141; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14214 = 10'h378 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11142; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14215 = 10'h379 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11143; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14216 = 10'h37a == _dirty_T_1 ? _cache_data_T_13 : _GEN_11144; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14217 = 10'h37b == _dirty_T_1 ? _cache_data_T_13 : _GEN_11145; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14218 = 10'h37c == _dirty_T_1 ? _cache_data_T_13 : _GEN_11146; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14219 = 10'h37d == _dirty_T_1 ? _cache_data_T_13 : _GEN_11147; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14220 = 10'h37e == _dirty_T_1 ? _cache_data_T_13 : _GEN_11148; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14221 = 10'h37f == _dirty_T_1 ? _cache_data_T_13 : _GEN_11149; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14222 = 10'h380 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11150; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14223 = 10'h381 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11151; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14224 = 10'h382 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11152; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14225 = 10'h383 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11153; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14226 = 10'h384 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11154; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14227 = 10'h385 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11155; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14228 = 10'h386 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11156; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14229 = 10'h387 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11157; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14230 = 10'h388 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11158; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14231 = 10'h389 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11159; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14232 = 10'h38a == _dirty_T_1 ? _cache_data_T_13 : _GEN_11160; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14233 = 10'h38b == _dirty_T_1 ? _cache_data_T_13 : _GEN_11161; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14234 = 10'h38c == _dirty_T_1 ? _cache_data_T_13 : _GEN_11162; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14235 = 10'h38d == _dirty_T_1 ? _cache_data_T_13 : _GEN_11163; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14236 = 10'h38e == _dirty_T_1 ? _cache_data_T_13 : _GEN_11164; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14237 = 10'h38f == _dirty_T_1 ? _cache_data_T_13 : _GEN_11165; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14238 = 10'h390 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11166; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14239 = 10'h391 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11167; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14240 = 10'h392 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11168; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14241 = 10'h393 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11169; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14242 = 10'h394 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11170; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14243 = 10'h395 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11171; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14244 = 10'h396 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11172; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14245 = 10'h397 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11173; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14246 = 10'h398 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11174; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14247 = 10'h399 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11175; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14248 = 10'h39a == _dirty_T_1 ? _cache_data_T_13 : _GEN_11176; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14249 = 10'h39b == _dirty_T_1 ? _cache_data_T_13 : _GEN_11177; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14250 = 10'h39c == _dirty_T_1 ? _cache_data_T_13 : _GEN_11178; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14251 = 10'h39d == _dirty_T_1 ? _cache_data_T_13 : _GEN_11179; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14252 = 10'h39e == _dirty_T_1 ? _cache_data_T_13 : _GEN_11180; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14253 = 10'h39f == _dirty_T_1 ? _cache_data_T_13 : _GEN_11181; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14254 = 10'h3a0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11182; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14255 = 10'h3a1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11183; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14256 = 10'h3a2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11184; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14257 = 10'h3a3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11185; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14258 = 10'h3a4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11186; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14259 = 10'h3a5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11187; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14260 = 10'h3a6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11188; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14261 = 10'h3a7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11189; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14262 = 10'h3a8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11190; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14263 = 10'h3a9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11191; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14264 = 10'h3aa == _dirty_T_1 ? _cache_data_T_13 : _GEN_11192; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14265 = 10'h3ab == _dirty_T_1 ? _cache_data_T_13 : _GEN_11193; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14266 = 10'h3ac == _dirty_T_1 ? _cache_data_T_13 : _GEN_11194; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14267 = 10'h3ad == _dirty_T_1 ? _cache_data_T_13 : _GEN_11195; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14268 = 10'h3ae == _dirty_T_1 ? _cache_data_T_13 : _GEN_11196; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14269 = 10'h3af == _dirty_T_1 ? _cache_data_T_13 : _GEN_11197; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14270 = 10'h3b0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11198; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14271 = 10'h3b1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11199; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14272 = 10'h3b2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11200; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14273 = 10'h3b3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11201; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14274 = 10'h3b4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11202; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14275 = 10'h3b5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11203; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14276 = 10'h3b6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11204; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14277 = 10'h3b7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11205; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14278 = 10'h3b8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11206; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14279 = 10'h3b9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11207; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14280 = 10'h3ba == _dirty_T_1 ? _cache_data_T_13 : _GEN_11208; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14281 = 10'h3bb == _dirty_T_1 ? _cache_data_T_13 : _GEN_11209; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14282 = 10'h3bc == _dirty_T_1 ? _cache_data_T_13 : _GEN_11210; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14283 = 10'h3bd == _dirty_T_1 ? _cache_data_T_13 : _GEN_11211; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14284 = 10'h3be == _dirty_T_1 ? _cache_data_T_13 : _GEN_11212; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14285 = 10'h3bf == _dirty_T_1 ? _cache_data_T_13 : _GEN_11213; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14286 = 10'h3c0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11214; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14287 = 10'h3c1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11215; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14288 = 10'h3c2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11216; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14289 = 10'h3c3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11217; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14290 = 10'h3c4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11218; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14291 = 10'h3c5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11219; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14292 = 10'h3c6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11220; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14293 = 10'h3c7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11221; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14294 = 10'h3c8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11222; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14295 = 10'h3c9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11223; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14296 = 10'h3ca == _dirty_T_1 ? _cache_data_T_13 : _GEN_11224; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14297 = 10'h3cb == _dirty_T_1 ? _cache_data_T_13 : _GEN_11225; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14298 = 10'h3cc == _dirty_T_1 ? _cache_data_T_13 : _GEN_11226; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14299 = 10'h3cd == _dirty_T_1 ? _cache_data_T_13 : _GEN_11227; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14300 = 10'h3ce == _dirty_T_1 ? _cache_data_T_13 : _GEN_11228; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14301 = 10'h3cf == _dirty_T_1 ? _cache_data_T_13 : _GEN_11229; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14302 = 10'h3d0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11230; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14303 = 10'h3d1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11231; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14304 = 10'h3d2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11232; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14305 = 10'h3d3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11233; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14306 = 10'h3d4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11234; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14307 = 10'h3d5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11235; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14308 = 10'h3d6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11236; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14309 = 10'h3d7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11237; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14310 = 10'h3d8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11238; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14311 = 10'h3d9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11239; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14312 = 10'h3da == _dirty_T_1 ? _cache_data_T_13 : _GEN_11240; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14313 = 10'h3db == _dirty_T_1 ? _cache_data_T_13 : _GEN_11241; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14314 = 10'h3dc == _dirty_T_1 ? _cache_data_T_13 : _GEN_11242; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14315 = 10'h3dd == _dirty_T_1 ? _cache_data_T_13 : _GEN_11243; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14316 = 10'h3de == _dirty_T_1 ? _cache_data_T_13 : _GEN_11244; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14317 = 10'h3df == _dirty_T_1 ? _cache_data_T_13 : _GEN_11245; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14318 = 10'h3e0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11246; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14319 = 10'h3e1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11247; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14320 = 10'h3e2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11248; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14321 = 10'h3e3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11249; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14322 = 10'h3e4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11250; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14323 = 10'h3e5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11251; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14324 = 10'h3e6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11252; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14325 = 10'h3e7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11253; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14326 = 10'h3e8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11254; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14327 = 10'h3e9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11255; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14328 = 10'h3ea == _dirty_T_1 ? _cache_data_T_13 : _GEN_11256; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14329 = 10'h3eb == _dirty_T_1 ? _cache_data_T_13 : _GEN_11257; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14330 = 10'h3ec == _dirty_T_1 ? _cache_data_T_13 : _GEN_11258; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14331 = 10'h3ed == _dirty_T_1 ? _cache_data_T_13 : _GEN_11259; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14332 = 10'h3ee == _dirty_T_1 ? _cache_data_T_13 : _GEN_11260; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14333 = 10'h3ef == _dirty_T_1 ? _cache_data_T_13 : _GEN_11261; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14334 = 10'h3f0 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11262; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14335 = 10'h3f1 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11263; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14336 = 10'h3f2 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11264; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14337 = 10'h3f3 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11265; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14338 = 10'h3f4 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11266; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14339 = 10'h3f5 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11267; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14340 = 10'h3f6 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11268; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14341 = 10'h3f7 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11269; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14342 = 10'h3f8 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11270; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14343 = 10'h3f9 == _dirty_T_1 ? _cache_data_T_13 : _GEN_11271; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14344 = 10'h3fa == _dirty_T_1 ? _cache_data_T_13 : _GEN_11272; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14345 = 10'h3fb == _dirty_T_1 ? _cache_data_T_13 : _GEN_11273; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14346 = 10'h3fc == _dirty_T_1 ? _cache_data_T_13 : _GEN_11274; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14347 = 10'h3fd == _dirty_T_1 ? _cache_data_T_13 : _GEN_11275; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14348 = 10'h3fe == _dirty_T_1 ? _cache_data_T_13 : _GEN_11276; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14349 = 10'h3ff == _dirty_T_1 ? _cache_data_T_13 : _GEN_11277; // @[icache.scala 139:{33,33}]
  wire [184:0] _GEN_14350 = lookup & dirty ? _GEN_13326 : _GEN_10254; // @[icache.scala 138:25]
  wire [184:0] _GEN_14351 = lookup & dirty ? _GEN_13327 : _GEN_10255; // @[icache.scala 138:25]
  wire [184:0] _GEN_14352 = lookup & dirty ? _GEN_13328 : _GEN_10256; // @[icache.scala 138:25]
  wire [184:0] _GEN_14353 = lookup & dirty ? _GEN_13329 : _GEN_10257; // @[icache.scala 138:25]
  wire [184:0] _GEN_14354 = lookup & dirty ? _GEN_13330 : _GEN_10258; // @[icache.scala 138:25]
  wire [184:0] _GEN_14355 = lookup & dirty ? _GEN_13331 : _GEN_10259; // @[icache.scala 138:25]
  wire [184:0] _GEN_14356 = lookup & dirty ? _GEN_13332 : _GEN_10260; // @[icache.scala 138:25]
  wire [184:0] _GEN_14357 = lookup & dirty ? _GEN_13333 : _GEN_10261; // @[icache.scala 138:25]
  wire [184:0] _GEN_14358 = lookup & dirty ? _GEN_13334 : _GEN_10262; // @[icache.scala 138:25]
  wire [184:0] _GEN_14359 = lookup & dirty ? _GEN_13335 : _GEN_10263; // @[icache.scala 138:25]
  wire [184:0] _GEN_14360 = lookup & dirty ? _GEN_13336 : _GEN_10264; // @[icache.scala 138:25]
  wire [184:0] _GEN_14361 = lookup & dirty ? _GEN_13337 : _GEN_10265; // @[icache.scala 138:25]
  wire [184:0] _GEN_14362 = lookup & dirty ? _GEN_13338 : _GEN_10266; // @[icache.scala 138:25]
  wire [184:0] _GEN_14363 = lookup & dirty ? _GEN_13339 : _GEN_10267; // @[icache.scala 138:25]
  wire [184:0] _GEN_14364 = lookup & dirty ? _GEN_13340 : _GEN_10268; // @[icache.scala 138:25]
  wire [184:0] _GEN_14365 = lookup & dirty ? _GEN_13341 : _GEN_10269; // @[icache.scala 138:25]
  wire [184:0] _GEN_14366 = lookup & dirty ? _GEN_13342 : _GEN_10270; // @[icache.scala 138:25]
  wire [184:0] _GEN_14367 = lookup & dirty ? _GEN_13343 : _GEN_10271; // @[icache.scala 138:25]
  wire [184:0] _GEN_14368 = lookup & dirty ? _GEN_13344 : _GEN_10272; // @[icache.scala 138:25]
  wire [184:0] _GEN_14369 = lookup & dirty ? _GEN_13345 : _GEN_10273; // @[icache.scala 138:25]
  wire [184:0] _GEN_14370 = lookup & dirty ? _GEN_13346 : _GEN_10274; // @[icache.scala 138:25]
  wire [184:0] _GEN_14371 = lookup & dirty ? _GEN_13347 : _GEN_10275; // @[icache.scala 138:25]
  wire [184:0] _GEN_14372 = lookup & dirty ? _GEN_13348 : _GEN_10276; // @[icache.scala 138:25]
  wire [184:0] _GEN_14373 = lookup & dirty ? _GEN_13349 : _GEN_10277; // @[icache.scala 138:25]
  wire [184:0] _GEN_14374 = lookup & dirty ? _GEN_13350 : _GEN_10278; // @[icache.scala 138:25]
  wire [184:0] _GEN_14375 = lookup & dirty ? _GEN_13351 : _GEN_10279; // @[icache.scala 138:25]
  wire [184:0] _GEN_14376 = lookup & dirty ? _GEN_13352 : _GEN_10280; // @[icache.scala 138:25]
  wire [184:0] _GEN_14377 = lookup & dirty ? _GEN_13353 : _GEN_10281; // @[icache.scala 138:25]
  wire [184:0] _GEN_14378 = lookup & dirty ? _GEN_13354 : _GEN_10282; // @[icache.scala 138:25]
  wire [184:0] _GEN_14379 = lookup & dirty ? _GEN_13355 : _GEN_10283; // @[icache.scala 138:25]
  wire [184:0] _GEN_14380 = lookup & dirty ? _GEN_13356 : _GEN_10284; // @[icache.scala 138:25]
  wire [184:0] _GEN_14381 = lookup & dirty ? _GEN_13357 : _GEN_10285; // @[icache.scala 138:25]
  wire [184:0] _GEN_14382 = lookup & dirty ? _GEN_13358 : _GEN_10286; // @[icache.scala 138:25]
  wire [184:0] _GEN_14383 = lookup & dirty ? _GEN_13359 : _GEN_10287; // @[icache.scala 138:25]
  wire [184:0] _GEN_14384 = lookup & dirty ? _GEN_13360 : _GEN_10288; // @[icache.scala 138:25]
  wire [184:0] _GEN_14385 = lookup & dirty ? _GEN_13361 : _GEN_10289; // @[icache.scala 138:25]
  wire [184:0] _GEN_14386 = lookup & dirty ? _GEN_13362 : _GEN_10290; // @[icache.scala 138:25]
  wire [184:0] _GEN_14387 = lookup & dirty ? _GEN_13363 : _GEN_10291; // @[icache.scala 138:25]
  wire [184:0] _GEN_14388 = lookup & dirty ? _GEN_13364 : _GEN_10292; // @[icache.scala 138:25]
  wire [184:0] _GEN_14389 = lookup & dirty ? _GEN_13365 : _GEN_10293; // @[icache.scala 138:25]
  wire [184:0] _GEN_14390 = lookup & dirty ? _GEN_13366 : _GEN_10294; // @[icache.scala 138:25]
  wire [184:0] _GEN_14391 = lookup & dirty ? _GEN_13367 : _GEN_10295; // @[icache.scala 138:25]
  wire [184:0] _GEN_14392 = lookup & dirty ? _GEN_13368 : _GEN_10296; // @[icache.scala 138:25]
  wire [184:0] _GEN_14393 = lookup & dirty ? _GEN_13369 : _GEN_10297; // @[icache.scala 138:25]
  wire [184:0] _GEN_14394 = lookup & dirty ? _GEN_13370 : _GEN_10298; // @[icache.scala 138:25]
  wire [184:0] _GEN_14395 = lookup & dirty ? _GEN_13371 : _GEN_10299; // @[icache.scala 138:25]
  wire [184:0] _GEN_14396 = lookup & dirty ? _GEN_13372 : _GEN_10300; // @[icache.scala 138:25]
  wire [184:0] _GEN_14397 = lookup & dirty ? _GEN_13373 : _GEN_10301; // @[icache.scala 138:25]
  wire [184:0] _GEN_14398 = lookup & dirty ? _GEN_13374 : _GEN_10302; // @[icache.scala 138:25]
  wire [184:0] _GEN_14399 = lookup & dirty ? _GEN_13375 : _GEN_10303; // @[icache.scala 138:25]
  wire [184:0] _GEN_14400 = lookup & dirty ? _GEN_13376 : _GEN_10304; // @[icache.scala 138:25]
  wire [184:0] _GEN_14401 = lookup & dirty ? _GEN_13377 : _GEN_10305; // @[icache.scala 138:25]
  wire [184:0] _GEN_14402 = lookup & dirty ? _GEN_13378 : _GEN_10306; // @[icache.scala 138:25]
  wire [184:0] _GEN_14403 = lookup & dirty ? _GEN_13379 : _GEN_10307; // @[icache.scala 138:25]
  wire [184:0] _GEN_14404 = lookup & dirty ? _GEN_13380 : _GEN_10308; // @[icache.scala 138:25]
  wire [184:0] _GEN_14405 = lookup & dirty ? _GEN_13381 : _GEN_10309; // @[icache.scala 138:25]
  wire [184:0] _GEN_14406 = lookup & dirty ? _GEN_13382 : _GEN_10310; // @[icache.scala 138:25]
  wire [184:0] _GEN_14407 = lookup & dirty ? _GEN_13383 : _GEN_10311; // @[icache.scala 138:25]
  wire [184:0] _GEN_14408 = lookup & dirty ? _GEN_13384 : _GEN_10312; // @[icache.scala 138:25]
  wire [184:0] _GEN_14409 = lookup & dirty ? _GEN_13385 : _GEN_10313; // @[icache.scala 138:25]
  wire [184:0] _GEN_14410 = lookup & dirty ? _GEN_13386 : _GEN_10314; // @[icache.scala 138:25]
  wire [184:0] _GEN_14411 = lookup & dirty ? _GEN_13387 : _GEN_10315; // @[icache.scala 138:25]
  wire [184:0] _GEN_14412 = lookup & dirty ? _GEN_13388 : _GEN_10316; // @[icache.scala 138:25]
  wire [184:0] _GEN_14413 = lookup & dirty ? _GEN_13389 : _GEN_10317; // @[icache.scala 138:25]
  wire [184:0] _GEN_14414 = lookup & dirty ? _GEN_13390 : _GEN_10318; // @[icache.scala 138:25]
  wire [184:0] _GEN_14415 = lookup & dirty ? _GEN_13391 : _GEN_10319; // @[icache.scala 138:25]
  wire [184:0] _GEN_14416 = lookup & dirty ? _GEN_13392 : _GEN_10320; // @[icache.scala 138:25]
  wire [184:0] _GEN_14417 = lookup & dirty ? _GEN_13393 : _GEN_10321; // @[icache.scala 138:25]
  wire [184:0] _GEN_14418 = lookup & dirty ? _GEN_13394 : _GEN_10322; // @[icache.scala 138:25]
  wire [184:0] _GEN_14419 = lookup & dirty ? _GEN_13395 : _GEN_10323; // @[icache.scala 138:25]
  wire [184:0] _GEN_14420 = lookup & dirty ? _GEN_13396 : _GEN_10324; // @[icache.scala 138:25]
  wire [184:0] _GEN_14421 = lookup & dirty ? _GEN_13397 : _GEN_10325; // @[icache.scala 138:25]
  wire [184:0] _GEN_14422 = lookup & dirty ? _GEN_13398 : _GEN_10326; // @[icache.scala 138:25]
  wire [184:0] _GEN_14423 = lookup & dirty ? _GEN_13399 : _GEN_10327; // @[icache.scala 138:25]
  wire [184:0] _GEN_14424 = lookup & dirty ? _GEN_13400 : _GEN_10328; // @[icache.scala 138:25]
  wire [184:0] _GEN_14425 = lookup & dirty ? _GEN_13401 : _GEN_10329; // @[icache.scala 138:25]
  wire [184:0] _GEN_14426 = lookup & dirty ? _GEN_13402 : _GEN_10330; // @[icache.scala 138:25]
  wire [184:0] _GEN_14427 = lookup & dirty ? _GEN_13403 : _GEN_10331; // @[icache.scala 138:25]
  wire [184:0] _GEN_14428 = lookup & dirty ? _GEN_13404 : _GEN_10332; // @[icache.scala 138:25]
  wire [184:0] _GEN_14429 = lookup & dirty ? _GEN_13405 : _GEN_10333; // @[icache.scala 138:25]
  wire [184:0] _GEN_14430 = lookup & dirty ? _GEN_13406 : _GEN_10334; // @[icache.scala 138:25]
  wire [184:0] _GEN_14431 = lookup & dirty ? _GEN_13407 : _GEN_10335; // @[icache.scala 138:25]
  wire [184:0] _GEN_14432 = lookup & dirty ? _GEN_13408 : _GEN_10336; // @[icache.scala 138:25]
  wire [184:0] _GEN_14433 = lookup & dirty ? _GEN_13409 : _GEN_10337; // @[icache.scala 138:25]
  wire [184:0] _GEN_14434 = lookup & dirty ? _GEN_13410 : _GEN_10338; // @[icache.scala 138:25]
  wire [184:0] _GEN_14435 = lookup & dirty ? _GEN_13411 : _GEN_10339; // @[icache.scala 138:25]
  wire [184:0] _GEN_14436 = lookup & dirty ? _GEN_13412 : _GEN_10340; // @[icache.scala 138:25]
  wire [184:0] _GEN_14437 = lookup & dirty ? _GEN_13413 : _GEN_10341; // @[icache.scala 138:25]
  wire [184:0] _GEN_14438 = lookup & dirty ? _GEN_13414 : _GEN_10342; // @[icache.scala 138:25]
  wire [184:0] _GEN_14439 = lookup & dirty ? _GEN_13415 : _GEN_10343; // @[icache.scala 138:25]
  wire [184:0] _GEN_14440 = lookup & dirty ? _GEN_13416 : _GEN_10344; // @[icache.scala 138:25]
  wire [184:0] _GEN_14441 = lookup & dirty ? _GEN_13417 : _GEN_10345; // @[icache.scala 138:25]
  wire [184:0] _GEN_14442 = lookup & dirty ? _GEN_13418 : _GEN_10346; // @[icache.scala 138:25]
  wire [184:0] _GEN_14443 = lookup & dirty ? _GEN_13419 : _GEN_10347; // @[icache.scala 138:25]
  wire [184:0] _GEN_14444 = lookup & dirty ? _GEN_13420 : _GEN_10348; // @[icache.scala 138:25]
  wire [184:0] _GEN_14445 = lookup & dirty ? _GEN_13421 : _GEN_10349; // @[icache.scala 138:25]
  wire [184:0] _GEN_14446 = lookup & dirty ? _GEN_13422 : _GEN_10350; // @[icache.scala 138:25]
  wire [184:0] _GEN_14447 = lookup & dirty ? _GEN_13423 : _GEN_10351; // @[icache.scala 138:25]
  wire [184:0] _GEN_14448 = lookup & dirty ? _GEN_13424 : _GEN_10352; // @[icache.scala 138:25]
  wire [184:0] _GEN_14449 = lookup & dirty ? _GEN_13425 : _GEN_10353; // @[icache.scala 138:25]
  wire [184:0] _GEN_14450 = lookup & dirty ? _GEN_13426 : _GEN_10354; // @[icache.scala 138:25]
  wire [184:0] _GEN_14451 = lookup & dirty ? _GEN_13427 : _GEN_10355; // @[icache.scala 138:25]
  wire [184:0] _GEN_14452 = lookup & dirty ? _GEN_13428 : _GEN_10356; // @[icache.scala 138:25]
  wire [184:0] _GEN_14453 = lookup & dirty ? _GEN_13429 : _GEN_10357; // @[icache.scala 138:25]
  wire [184:0] _GEN_14454 = lookup & dirty ? _GEN_13430 : _GEN_10358; // @[icache.scala 138:25]
  wire [184:0] _GEN_14455 = lookup & dirty ? _GEN_13431 : _GEN_10359; // @[icache.scala 138:25]
  wire [184:0] _GEN_14456 = lookup & dirty ? _GEN_13432 : _GEN_10360; // @[icache.scala 138:25]
  wire [184:0] _GEN_14457 = lookup & dirty ? _GEN_13433 : _GEN_10361; // @[icache.scala 138:25]
  wire [184:0] _GEN_14458 = lookup & dirty ? _GEN_13434 : _GEN_10362; // @[icache.scala 138:25]
  wire [184:0] _GEN_14459 = lookup & dirty ? _GEN_13435 : _GEN_10363; // @[icache.scala 138:25]
  wire [184:0] _GEN_14460 = lookup & dirty ? _GEN_13436 : _GEN_10364; // @[icache.scala 138:25]
  wire [184:0] _GEN_14461 = lookup & dirty ? _GEN_13437 : _GEN_10365; // @[icache.scala 138:25]
  wire [184:0] _GEN_14462 = lookup & dirty ? _GEN_13438 : _GEN_10366; // @[icache.scala 138:25]
  wire [184:0] _GEN_14463 = lookup & dirty ? _GEN_13439 : _GEN_10367; // @[icache.scala 138:25]
  wire [184:0] _GEN_14464 = lookup & dirty ? _GEN_13440 : _GEN_10368; // @[icache.scala 138:25]
  wire [184:0] _GEN_14465 = lookup & dirty ? _GEN_13441 : _GEN_10369; // @[icache.scala 138:25]
  wire [184:0] _GEN_14466 = lookup & dirty ? _GEN_13442 : _GEN_10370; // @[icache.scala 138:25]
  wire [184:0] _GEN_14467 = lookup & dirty ? _GEN_13443 : _GEN_10371; // @[icache.scala 138:25]
  wire [184:0] _GEN_14468 = lookup & dirty ? _GEN_13444 : _GEN_10372; // @[icache.scala 138:25]
  wire [184:0] _GEN_14469 = lookup & dirty ? _GEN_13445 : _GEN_10373; // @[icache.scala 138:25]
  wire [184:0] _GEN_14470 = lookup & dirty ? _GEN_13446 : _GEN_10374; // @[icache.scala 138:25]
  wire [184:0] _GEN_14471 = lookup & dirty ? _GEN_13447 : _GEN_10375; // @[icache.scala 138:25]
  wire [184:0] _GEN_14472 = lookup & dirty ? _GEN_13448 : _GEN_10376; // @[icache.scala 138:25]
  wire [184:0] _GEN_14473 = lookup & dirty ? _GEN_13449 : _GEN_10377; // @[icache.scala 138:25]
  wire [184:0] _GEN_14474 = lookup & dirty ? _GEN_13450 : _GEN_10378; // @[icache.scala 138:25]
  wire [184:0] _GEN_14475 = lookup & dirty ? _GEN_13451 : _GEN_10379; // @[icache.scala 138:25]
  wire [184:0] _GEN_14476 = lookup & dirty ? _GEN_13452 : _GEN_10380; // @[icache.scala 138:25]
  wire [184:0] _GEN_14477 = lookup & dirty ? _GEN_13453 : _GEN_10381; // @[icache.scala 138:25]
  wire [184:0] _GEN_14478 = lookup & dirty ? _GEN_13454 : _GEN_10382; // @[icache.scala 138:25]
  wire [184:0] _GEN_14479 = lookup & dirty ? _GEN_13455 : _GEN_10383; // @[icache.scala 138:25]
  wire [184:0] _GEN_14480 = lookup & dirty ? _GEN_13456 : _GEN_10384; // @[icache.scala 138:25]
  wire [184:0] _GEN_14481 = lookup & dirty ? _GEN_13457 : _GEN_10385; // @[icache.scala 138:25]
  wire [184:0] _GEN_14482 = lookup & dirty ? _GEN_13458 : _GEN_10386; // @[icache.scala 138:25]
  wire [184:0] _GEN_14483 = lookup & dirty ? _GEN_13459 : _GEN_10387; // @[icache.scala 138:25]
  wire [184:0] _GEN_14484 = lookup & dirty ? _GEN_13460 : _GEN_10388; // @[icache.scala 138:25]
  wire [184:0] _GEN_14485 = lookup & dirty ? _GEN_13461 : _GEN_10389; // @[icache.scala 138:25]
  wire [184:0] _GEN_14486 = lookup & dirty ? _GEN_13462 : _GEN_10390; // @[icache.scala 138:25]
  wire [184:0] _GEN_14487 = lookup & dirty ? _GEN_13463 : _GEN_10391; // @[icache.scala 138:25]
  wire [184:0] _GEN_14488 = lookup & dirty ? _GEN_13464 : _GEN_10392; // @[icache.scala 138:25]
  wire [184:0] _GEN_14489 = lookup & dirty ? _GEN_13465 : _GEN_10393; // @[icache.scala 138:25]
  wire [184:0] _GEN_14490 = lookup & dirty ? _GEN_13466 : _GEN_10394; // @[icache.scala 138:25]
  wire [184:0] _GEN_14491 = lookup & dirty ? _GEN_13467 : _GEN_10395; // @[icache.scala 138:25]
  wire [184:0] _GEN_14492 = lookup & dirty ? _GEN_13468 : _GEN_10396; // @[icache.scala 138:25]
  wire [184:0] _GEN_14493 = lookup & dirty ? _GEN_13469 : _GEN_10397; // @[icache.scala 138:25]
  wire [184:0] _GEN_14494 = lookup & dirty ? _GEN_13470 : _GEN_10398; // @[icache.scala 138:25]
  wire [184:0] _GEN_14495 = lookup & dirty ? _GEN_13471 : _GEN_10399; // @[icache.scala 138:25]
  wire [184:0] _GEN_14496 = lookup & dirty ? _GEN_13472 : _GEN_10400; // @[icache.scala 138:25]
  wire [184:0] _GEN_14497 = lookup & dirty ? _GEN_13473 : _GEN_10401; // @[icache.scala 138:25]
  wire [184:0] _GEN_14498 = lookup & dirty ? _GEN_13474 : _GEN_10402; // @[icache.scala 138:25]
  wire [184:0] _GEN_14499 = lookup & dirty ? _GEN_13475 : _GEN_10403; // @[icache.scala 138:25]
  wire [184:0] _GEN_14500 = lookup & dirty ? _GEN_13476 : _GEN_10404; // @[icache.scala 138:25]
  wire [184:0] _GEN_14501 = lookup & dirty ? _GEN_13477 : _GEN_10405; // @[icache.scala 138:25]
  wire [184:0] _GEN_14502 = lookup & dirty ? _GEN_13478 : _GEN_10406; // @[icache.scala 138:25]
  wire [184:0] _GEN_14503 = lookup & dirty ? _GEN_13479 : _GEN_10407; // @[icache.scala 138:25]
  wire [184:0] _GEN_14504 = lookup & dirty ? _GEN_13480 : _GEN_10408; // @[icache.scala 138:25]
  wire [184:0] _GEN_14505 = lookup & dirty ? _GEN_13481 : _GEN_10409; // @[icache.scala 138:25]
  wire [184:0] _GEN_14506 = lookup & dirty ? _GEN_13482 : _GEN_10410; // @[icache.scala 138:25]
  wire [184:0] _GEN_14507 = lookup & dirty ? _GEN_13483 : _GEN_10411; // @[icache.scala 138:25]
  wire [184:0] _GEN_14508 = lookup & dirty ? _GEN_13484 : _GEN_10412; // @[icache.scala 138:25]
  wire [184:0] _GEN_14509 = lookup & dirty ? _GEN_13485 : _GEN_10413; // @[icache.scala 138:25]
  wire [184:0] _GEN_14510 = lookup & dirty ? _GEN_13486 : _GEN_10414; // @[icache.scala 138:25]
  wire [184:0] _GEN_14511 = lookup & dirty ? _GEN_13487 : _GEN_10415; // @[icache.scala 138:25]
  wire [184:0] _GEN_14512 = lookup & dirty ? _GEN_13488 : _GEN_10416; // @[icache.scala 138:25]
  wire [184:0] _GEN_14513 = lookup & dirty ? _GEN_13489 : _GEN_10417; // @[icache.scala 138:25]
  wire [184:0] _GEN_14514 = lookup & dirty ? _GEN_13490 : _GEN_10418; // @[icache.scala 138:25]
  wire [184:0] _GEN_14515 = lookup & dirty ? _GEN_13491 : _GEN_10419; // @[icache.scala 138:25]
  wire [184:0] _GEN_14516 = lookup & dirty ? _GEN_13492 : _GEN_10420; // @[icache.scala 138:25]
  wire [184:0] _GEN_14517 = lookup & dirty ? _GEN_13493 : _GEN_10421; // @[icache.scala 138:25]
  wire [184:0] _GEN_14518 = lookup & dirty ? _GEN_13494 : _GEN_10422; // @[icache.scala 138:25]
  wire [184:0] _GEN_14519 = lookup & dirty ? _GEN_13495 : _GEN_10423; // @[icache.scala 138:25]
  wire [184:0] _GEN_14520 = lookup & dirty ? _GEN_13496 : _GEN_10424; // @[icache.scala 138:25]
  wire [184:0] _GEN_14521 = lookup & dirty ? _GEN_13497 : _GEN_10425; // @[icache.scala 138:25]
  wire [184:0] _GEN_14522 = lookup & dirty ? _GEN_13498 : _GEN_10426; // @[icache.scala 138:25]
  wire [184:0] _GEN_14523 = lookup & dirty ? _GEN_13499 : _GEN_10427; // @[icache.scala 138:25]
  wire [184:0] _GEN_14524 = lookup & dirty ? _GEN_13500 : _GEN_10428; // @[icache.scala 138:25]
  wire [184:0] _GEN_14525 = lookup & dirty ? _GEN_13501 : _GEN_10429; // @[icache.scala 138:25]
  wire [184:0] _GEN_14526 = lookup & dirty ? _GEN_13502 : _GEN_10430; // @[icache.scala 138:25]
  wire [184:0] _GEN_14527 = lookup & dirty ? _GEN_13503 : _GEN_10431; // @[icache.scala 138:25]
  wire [184:0] _GEN_14528 = lookup & dirty ? _GEN_13504 : _GEN_10432; // @[icache.scala 138:25]
  wire [184:0] _GEN_14529 = lookup & dirty ? _GEN_13505 : _GEN_10433; // @[icache.scala 138:25]
  wire [184:0] _GEN_14530 = lookup & dirty ? _GEN_13506 : _GEN_10434; // @[icache.scala 138:25]
  wire [184:0] _GEN_14531 = lookup & dirty ? _GEN_13507 : _GEN_10435; // @[icache.scala 138:25]
  wire [184:0] _GEN_14532 = lookup & dirty ? _GEN_13508 : _GEN_10436; // @[icache.scala 138:25]
  wire [184:0] _GEN_14533 = lookup & dirty ? _GEN_13509 : _GEN_10437; // @[icache.scala 138:25]
  wire [184:0] _GEN_14534 = lookup & dirty ? _GEN_13510 : _GEN_10438; // @[icache.scala 138:25]
  wire [184:0] _GEN_14535 = lookup & dirty ? _GEN_13511 : _GEN_10439; // @[icache.scala 138:25]
  wire [184:0] _GEN_14536 = lookup & dirty ? _GEN_13512 : _GEN_10440; // @[icache.scala 138:25]
  wire [184:0] _GEN_14537 = lookup & dirty ? _GEN_13513 : _GEN_10441; // @[icache.scala 138:25]
  wire [184:0] _GEN_14538 = lookup & dirty ? _GEN_13514 : _GEN_10442; // @[icache.scala 138:25]
  wire [184:0] _GEN_14539 = lookup & dirty ? _GEN_13515 : _GEN_10443; // @[icache.scala 138:25]
  wire [184:0] _GEN_14540 = lookup & dirty ? _GEN_13516 : _GEN_10444; // @[icache.scala 138:25]
  wire [184:0] _GEN_14541 = lookup & dirty ? _GEN_13517 : _GEN_10445; // @[icache.scala 138:25]
  wire [184:0] _GEN_14542 = lookup & dirty ? _GEN_13518 : _GEN_10446; // @[icache.scala 138:25]
  wire [184:0] _GEN_14543 = lookup & dirty ? _GEN_13519 : _GEN_10447; // @[icache.scala 138:25]
  wire [184:0] _GEN_14544 = lookup & dirty ? _GEN_13520 : _GEN_10448; // @[icache.scala 138:25]
  wire [184:0] _GEN_14545 = lookup & dirty ? _GEN_13521 : _GEN_10449; // @[icache.scala 138:25]
  wire [184:0] _GEN_14546 = lookup & dirty ? _GEN_13522 : _GEN_10450; // @[icache.scala 138:25]
  wire [184:0] _GEN_14547 = lookup & dirty ? _GEN_13523 : _GEN_10451; // @[icache.scala 138:25]
  wire [184:0] _GEN_14548 = lookup & dirty ? _GEN_13524 : _GEN_10452; // @[icache.scala 138:25]
  wire [184:0] _GEN_14549 = lookup & dirty ? _GEN_13525 : _GEN_10453; // @[icache.scala 138:25]
  wire [184:0] _GEN_14550 = lookup & dirty ? _GEN_13526 : _GEN_10454; // @[icache.scala 138:25]
  wire [184:0] _GEN_14551 = lookup & dirty ? _GEN_13527 : _GEN_10455; // @[icache.scala 138:25]
  wire [184:0] _GEN_14552 = lookup & dirty ? _GEN_13528 : _GEN_10456; // @[icache.scala 138:25]
  wire [184:0] _GEN_14553 = lookup & dirty ? _GEN_13529 : _GEN_10457; // @[icache.scala 138:25]
  wire [184:0] _GEN_14554 = lookup & dirty ? _GEN_13530 : _GEN_10458; // @[icache.scala 138:25]
  wire [184:0] _GEN_14555 = lookup & dirty ? _GEN_13531 : _GEN_10459; // @[icache.scala 138:25]
  wire [184:0] _GEN_14556 = lookup & dirty ? _GEN_13532 : _GEN_10460; // @[icache.scala 138:25]
  wire [184:0] _GEN_14557 = lookup & dirty ? _GEN_13533 : _GEN_10461; // @[icache.scala 138:25]
  wire [184:0] _GEN_14558 = lookup & dirty ? _GEN_13534 : _GEN_10462; // @[icache.scala 138:25]
  wire [184:0] _GEN_14559 = lookup & dirty ? _GEN_13535 : _GEN_10463; // @[icache.scala 138:25]
  wire [184:0] _GEN_14560 = lookup & dirty ? _GEN_13536 : _GEN_10464; // @[icache.scala 138:25]
  wire [184:0] _GEN_14561 = lookup & dirty ? _GEN_13537 : _GEN_10465; // @[icache.scala 138:25]
  wire [184:0] _GEN_14562 = lookup & dirty ? _GEN_13538 : _GEN_10466; // @[icache.scala 138:25]
  wire [184:0] _GEN_14563 = lookup & dirty ? _GEN_13539 : _GEN_10467; // @[icache.scala 138:25]
  wire [184:0] _GEN_14564 = lookup & dirty ? _GEN_13540 : _GEN_10468; // @[icache.scala 138:25]
  wire [184:0] _GEN_14565 = lookup & dirty ? _GEN_13541 : _GEN_10469; // @[icache.scala 138:25]
  wire [184:0] _GEN_14566 = lookup & dirty ? _GEN_13542 : _GEN_10470; // @[icache.scala 138:25]
  wire [184:0] _GEN_14567 = lookup & dirty ? _GEN_13543 : _GEN_10471; // @[icache.scala 138:25]
  wire [184:0] _GEN_14568 = lookup & dirty ? _GEN_13544 : _GEN_10472; // @[icache.scala 138:25]
  wire [184:0] _GEN_14569 = lookup & dirty ? _GEN_13545 : _GEN_10473; // @[icache.scala 138:25]
  wire [184:0] _GEN_14570 = lookup & dirty ? _GEN_13546 : _GEN_10474; // @[icache.scala 138:25]
  wire [184:0] _GEN_14571 = lookup & dirty ? _GEN_13547 : _GEN_10475; // @[icache.scala 138:25]
  wire [184:0] _GEN_14572 = lookup & dirty ? _GEN_13548 : _GEN_10476; // @[icache.scala 138:25]
  wire [184:0] _GEN_14573 = lookup & dirty ? _GEN_13549 : _GEN_10477; // @[icache.scala 138:25]
  wire [184:0] _GEN_14574 = lookup & dirty ? _GEN_13550 : _GEN_10478; // @[icache.scala 138:25]
  wire [184:0] _GEN_14575 = lookup & dirty ? _GEN_13551 : _GEN_10479; // @[icache.scala 138:25]
  wire [184:0] _GEN_14576 = lookup & dirty ? _GEN_13552 : _GEN_10480; // @[icache.scala 138:25]
  wire [184:0] _GEN_14577 = lookup & dirty ? _GEN_13553 : _GEN_10481; // @[icache.scala 138:25]
  wire [184:0] _GEN_14578 = lookup & dirty ? _GEN_13554 : _GEN_10482; // @[icache.scala 138:25]
  wire [184:0] _GEN_14579 = lookup & dirty ? _GEN_13555 : _GEN_10483; // @[icache.scala 138:25]
  wire [184:0] _GEN_14580 = lookup & dirty ? _GEN_13556 : _GEN_10484; // @[icache.scala 138:25]
  wire [184:0] _GEN_14581 = lookup & dirty ? _GEN_13557 : _GEN_10485; // @[icache.scala 138:25]
  wire [184:0] _GEN_14582 = lookup & dirty ? _GEN_13558 : _GEN_10486; // @[icache.scala 138:25]
  wire [184:0] _GEN_14583 = lookup & dirty ? _GEN_13559 : _GEN_10487; // @[icache.scala 138:25]
  wire [184:0] _GEN_14584 = lookup & dirty ? _GEN_13560 : _GEN_10488; // @[icache.scala 138:25]
  wire [184:0] _GEN_14585 = lookup & dirty ? _GEN_13561 : _GEN_10489; // @[icache.scala 138:25]
  wire [184:0] _GEN_14586 = lookup & dirty ? _GEN_13562 : _GEN_10490; // @[icache.scala 138:25]
  wire [184:0] _GEN_14587 = lookup & dirty ? _GEN_13563 : _GEN_10491; // @[icache.scala 138:25]
  wire [184:0] _GEN_14588 = lookup & dirty ? _GEN_13564 : _GEN_10492; // @[icache.scala 138:25]
  wire [184:0] _GEN_14589 = lookup & dirty ? _GEN_13565 : _GEN_10493; // @[icache.scala 138:25]
  wire [184:0] _GEN_14590 = lookup & dirty ? _GEN_13566 : _GEN_10494; // @[icache.scala 138:25]
  wire [184:0] _GEN_14591 = lookup & dirty ? _GEN_13567 : _GEN_10495; // @[icache.scala 138:25]
  wire [184:0] _GEN_14592 = lookup & dirty ? _GEN_13568 : _GEN_10496; // @[icache.scala 138:25]
  wire [184:0] _GEN_14593 = lookup & dirty ? _GEN_13569 : _GEN_10497; // @[icache.scala 138:25]
  wire [184:0] _GEN_14594 = lookup & dirty ? _GEN_13570 : _GEN_10498; // @[icache.scala 138:25]
  wire [184:0] _GEN_14595 = lookup & dirty ? _GEN_13571 : _GEN_10499; // @[icache.scala 138:25]
  wire [184:0] _GEN_14596 = lookup & dirty ? _GEN_13572 : _GEN_10500; // @[icache.scala 138:25]
  wire [184:0] _GEN_14597 = lookup & dirty ? _GEN_13573 : _GEN_10501; // @[icache.scala 138:25]
  wire [184:0] _GEN_14598 = lookup & dirty ? _GEN_13574 : _GEN_10502; // @[icache.scala 138:25]
  wire [184:0] _GEN_14599 = lookup & dirty ? _GEN_13575 : _GEN_10503; // @[icache.scala 138:25]
  wire [184:0] _GEN_14600 = lookup & dirty ? _GEN_13576 : _GEN_10504; // @[icache.scala 138:25]
  wire [184:0] _GEN_14601 = lookup & dirty ? _GEN_13577 : _GEN_10505; // @[icache.scala 138:25]
  wire [184:0] _GEN_14602 = lookup & dirty ? _GEN_13578 : _GEN_10506; // @[icache.scala 138:25]
  wire [184:0] _GEN_14603 = lookup & dirty ? _GEN_13579 : _GEN_10507; // @[icache.scala 138:25]
  wire [184:0] _GEN_14604 = lookup & dirty ? _GEN_13580 : _GEN_10508; // @[icache.scala 138:25]
  wire [184:0] _GEN_14605 = lookup & dirty ? _GEN_13581 : _GEN_10509; // @[icache.scala 138:25]
  wire [184:0] _GEN_14606 = lookup & dirty ? _GEN_13582 : _GEN_10510; // @[icache.scala 138:25]
  wire [184:0] _GEN_14607 = lookup & dirty ? _GEN_13583 : _GEN_10511; // @[icache.scala 138:25]
  wire [184:0] _GEN_14608 = lookup & dirty ? _GEN_13584 : _GEN_10512; // @[icache.scala 138:25]
  wire [184:0] _GEN_14609 = lookup & dirty ? _GEN_13585 : _GEN_10513; // @[icache.scala 138:25]
  wire [184:0] _GEN_14610 = lookup & dirty ? _GEN_13586 : _GEN_10514; // @[icache.scala 138:25]
  wire [184:0] _GEN_14611 = lookup & dirty ? _GEN_13587 : _GEN_10515; // @[icache.scala 138:25]
  wire [184:0] _GEN_14612 = lookup & dirty ? _GEN_13588 : _GEN_10516; // @[icache.scala 138:25]
  wire [184:0] _GEN_14613 = lookup & dirty ? _GEN_13589 : _GEN_10517; // @[icache.scala 138:25]
  wire [184:0] _GEN_14614 = lookup & dirty ? _GEN_13590 : _GEN_10518; // @[icache.scala 138:25]
  wire [184:0] _GEN_14615 = lookup & dirty ? _GEN_13591 : _GEN_10519; // @[icache.scala 138:25]
  wire [184:0] _GEN_14616 = lookup & dirty ? _GEN_13592 : _GEN_10520; // @[icache.scala 138:25]
  wire [184:0] _GEN_14617 = lookup & dirty ? _GEN_13593 : _GEN_10521; // @[icache.scala 138:25]
  wire [184:0] _GEN_14618 = lookup & dirty ? _GEN_13594 : _GEN_10522; // @[icache.scala 138:25]
  wire [184:0] _GEN_14619 = lookup & dirty ? _GEN_13595 : _GEN_10523; // @[icache.scala 138:25]
  wire [184:0] _GEN_14620 = lookup & dirty ? _GEN_13596 : _GEN_10524; // @[icache.scala 138:25]
  wire [184:0] _GEN_14621 = lookup & dirty ? _GEN_13597 : _GEN_10525; // @[icache.scala 138:25]
  wire [184:0] _GEN_14622 = lookup & dirty ? _GEN_13598 : _GEN_10526; // @[icache.scala 138:25]
  wire [184:0] _GEN_14623 = lookup & dirty ? _GEN_13599 : _GEN_10527; // @[icache.scala 138:25]
  wire [184:0] _GEN_14624 = lookup & dirty ? _GEN_13600 : _GEN_10528; // @[icache.scala 138:25]
  wire [184:0] _GEN_14625 = lookup & dirty ? _GEN_13601 : _GEN_10529; // @[icache.scala 138:25]
  wire [184:0] _GEN_14626 = lookup & dirty ? _GEN_13602 : _GEN_10530; // @[icache.scala 138:25]
  wire [184:0] _GEN_14627 = lookup & dirty ? _GEN_13603 : _GEN_10531; // @[icache.scala 138:25]
  wire [184:0] _GEN_14628 = lookup & dirty ? _GEN_13604 : _GEN_10532; // @[icache.scala 138:25]
  wire [184:0] _GEN_14629 = lookup & dirty ? _GEN_13605 : _GEN_10533; // @[icache.scala 138:25]
  wire [184:0] _GEN_14630 = lookup & dirty ? _GEN_13606 : _GEN_10534; // @[icache.scala 138:25]
  wire [184:0] _GEN_14631 = lookup & dirty ? _GEN_13607 : _GEN_10535; // @[icache.scala 138:25]
  wire [184:0] _GEN_14632 = lookup & dirty ? _GEN_13608 : _GEN_10536; // @[icache.scala 138:25]
  wire [184:0] _GEN_14633 = lookup & dirty ? _GEN_13609 : _GEN_10537; // @[icache.scala 138:25]
  wire [184:0] _GEN_14634 = lookup & dirty ? _GEN_13610 : _GEN_10538; // @[icache.scala 138:25]
  wire [184:0] _GEN_14635 = lookup & dirty ? _GEN_13611 : _GEN_10539; // @[icache.scala 138:25]
  wire [184:0] _GEN_14636 = lookup & dirty ? _GEN_13612 : _GEN_10540; // @[icache.scala 138:25]
  wire [184:0] _GEN_14637 = lookup & dirty ? _GEN_13613 : _GEN_10541; // @[icache.scala 138:25]
  wire [184:0] _GEN_14638 = lookup & dirty ? _GEN_13614 : _GEN_10542; // @[icache.scala 138:25]
  wire [184:0] _GEN_14639 = lookup & dirty ? _GEN_13615 : _GEN_10543; // @[icache.scala 138:25]
  wire [184:0] _GEN_14640 = lookup & dirty ? _GEN_13616 : _GEN_10544; // @[icache.scala 138:25]
  wire [184:0] _GEN_14641 = lookup & dirty ? _GEN_13617 : _GEN_10545; // @[icache.scala 138:25]
  wire [184:0] _GEN_14642 = lookup & dirty ? _GEN_13618 : _GEN_10546; // @[icache.scala 138:25]
  wire [184:0] _GEN_14643 = lookup & dirty ? _GEN_13619 : _GEN_10547; // @[icache.scala 138:25]
  wire [184:0] _GEN_14644 = lookup & dirty ? _GEN_13620 : _GEN_10548; // @[icache.scala 138:25]
  wire [184:0] _GEN_14645 = lookup & dirty ? _GEN_13621 : _GEN_10549; // @[icache.scala 138:25]
  wire [184:0] _GEN_14646 = lookup & dirty ? _GEN_13622 : _GEN_10550; // @[icache.scala 138:25]
  wire [184:0] _GEN_14647 = lookup & dirty ? _GEN_13623 : _GEN_10551; // @[icache.scala 138:25]
  wire [184:0] _GEN_14648 = lookup & dirty ? _GEN_13624 : _GEN_10552; // @[icache.scala 138:25]
  wire [184:0] _GEN_14649 = lookup & dirty ? _GEN_13625 : _GEN_10553; // @[icache.scala 138:25]
  wire [184:0] _GEN_14650 = lookup & dirty ? _GEN_13626 : _GEN_10554; // @[icache.scala 138:25]
  wire [184:0] _GEN_14651 = lookup & dirty ? _GEN_13627 : _GEN_10555; // @[icache.scala 138:25]
  wire [184:0] _GEN_14652 = lookup & dirty ? _GEN_13628 : _GEN_10556; // @[icache.scala 138:25]
  wire [184:0] _GEN_14653 = lookup & dirty ? _GEN_13629 : _GEN_10557; // @[icache.scala 138:25]
  wire [184:0] _GEN_14654 = lookup & dirty ? _GEN_13630 : _GEN_10558; // @[icache.scala 138:25]
  wire [184:0] _GEN_14655 = lookup & dirty ? _GEN_13631 : _GEN_10559; // @[icache.scala 138:25]
  wire [184:0] _GEN_14656 = lookup & dirty ? _GEN_13632 : _GEN_10560; // @[icache.scala 138:25]
  wire [184:0] _GEN_14657 = lookup & dirty ? _GEN_13633 : _GEN_10561; // @[icache.scala 138:25]
  wire [184:0] _GEN_14658 = lookup & dirty ? _GEN_13634 : _GEN_10562; // @[icache.scala 138:25]
  wire [184:0] _GEN_14659 = lookup & dirty ? _GEN_13635 : _GEN_10563; // @[icache.scala 138:25]
  wire [184:0] _GEN_14660 = lookup & dirty ? _GEN_13636 : _GEN_10564; // @[icache.scala 138:25]
  wire [184:0] _GEN_14661 = lookup & dirty ? _GEN_13637 : _GEN_10565; // @[icache.scala 138:25]
  wire [184:0] _GEN_14662 = lookup & dirty ? _GEN_13638 : _GEN_10566; // @[icache.scala 138:25]
  wire [184:0] _GEN_14663 = lookup & dirty ? _GEN_13639 : _GEN_10567; // @[icache.scala 138:25]
  wire [184:0] _GEN_14664 = lookup & dirty ? _GEN_13640 : _GEN_10568; // @[icache.scala 138:25]
  wire [184:0] _GEN_14665 = lookup & dirty ? _GEN_13641 : _GEN_10569; // @[icache.scala 138:25]
  wire [184:0] _GEN_14666 = lookup & dirty ? _GEN_13642 : _GEN_10570; // @[icache.scala 138:25]
  wire [184:0] _GEN_14667 = lookup & dirty ? _GEN_13643 : _GEN_10571; // @[icache.scala 138:25]
  wire [184:0] _GEN_14668 = lookup & dirty ? _GEN_13644 : _GEN_10572; // @[icache.scala 138:25]
  wire [184:0] _GEN_14669 = lookup & dirty ? _GEN_13645 : _GEN_10573; // @[icache.scala 138:25]
  wire [184:0] _GEN_14670 = lookup & dirty ? _GEN_13646 : _GEN_10574; // @[icache.scala 138:25]
  wire [184:0] _GEN_14671 = lookup & dirty ? _GEN_13647 : _GEN_10575; // @[icache.scala 138:25]
  wire [184:0] _GEN_14672 = lookup & dirty ? _GEN_13648 : _GEN_10576; // @[icache.scala 138:25]
  wire [184:0] _GEN_14673 = lookup & dirty ? _GEN_13649 : _GEN_10577; // @[icache.scala 138:25]
  wire [184:0] _GEN_14674 = lookup & dirty ? _GEN_13650 : _GEN_10578; // @[icache.scala 138:25]
  wire [184:0] _GEN_14675 = lookup & dirty ? _GEN_13651 : _GEN_10579; // @[icache.scala 138:25]
  wire [184:0] _GEN_14676 = lookup & dirty ? _GEN_13652 : _GEN_10580; // @[icache.scala 138:25]
  wire [184:0] _GEN_14677 = lookup & dirty ? _GEN_13653 : _GEN_10581; // @[icache.scala 138:25]
  wire [184:0] _GEN_14678 = lookup & dirty ? _GEN_13654 : _GEN_10582; // @[icache.scala 138:25]
  wire [184:0] _GEN_14679 = lookup & dirty ? _GEN_13655 : _GEN_10583; // @[icache.scala 138:25]
  wire [184:0] _GEN_14680 = lookup & dirty ? _GEN_13656 : _GEN_10584; // @[icache.scala 138:25]
  wire [184:0] _GEN_14681 = lookup & dirty ? _GEN_13657 : _GEN_10585; // @[icache.scala 138:25]
  wire [184:0] _GEN_14682 = lookup & dirty ? _GEN_13658 : _GEN_10586; // @[icache.scala 138:25]
  wire [184:0] _GEN_14683 = lookup & dirty ? _GEN_13659 : _GEN_10587; // @[icache.scala 138:25]
  wire [184:0] _GEN_14684 = lookup & dirty ? _GEN_13660 : _GEN_10588; // @[icache.scala 138:25]
  wire [184:0] _GEN_14685 = lookup & dirty ? _GEN_13661 : _GEN_10589; // @[icache.scala 138:25]
  wire [184:0] _GEN_14686 = lookup & dirty ? _GEN_13662 : _GEN_10590; // @[icache.scala 138:25]
  wire [184:0] _GEN_14687 = lookup & dirty ? _GEN_13663 : _GEN_10591; // @[icache.scala 138:25]
  wire [184:0] _GEN_14688 = lookup & dirty ? _GEN_13664 : _GEN_10592; // @[icache.scala 138:25]
  wire [184:0] _GEN_14689 = lookup & dirty ? _GEN_13665 : _GEN_10593; // @[icache.scala 138:25]
  wire [184:0] _GEN_14690 = lookup & dirty ? _GEN_13666 : _GEN_10594; // @[icache.scala 138:25]
  wire [184:0] _GEN_14691 = lookup & dirty ? _GEN_13667 : _GEN_10595; // @[icache.scala 138:25]
  wire [184:0] _GEN_14692 = lookup & dirty ? _GEN_13668 : _GEN_10596; // @[icache.scala 138:25]
  wire [184:0] _GEN_14693 = lookup & dirty ? _GEN_13669 : _GEN_10597; // @[icache.scala 138:25]
  wire [184:0] _GEN_14694 = lookup & dirty ? _GEN_13670 : _GEN_10598; // @[icache.scala 138:25]
  wire [184:0] _GEN_14695 = lookup & dirty ? _GEN_13671 : _GEN_10599; // @[icache.scala 138:25]
  wire [184:0] _GEN_14696 = lookup & dirty ? _GEN_13672 : _GEN_10600; // @[icache.scala 138:25]
  wire [184:0] _GEN_14697 = lookup & dirty ? _GEN_13673 : _GEN_10601; // @[icache.scala 138:25]
  wire [184:0] _GEN_14698 = lookup & dirty ? _GEN_13674 : _GEN_10602; // @[icache.scala 138:25]
  wire [184:0] _GEN_14699 = lookup & dirty ? _GEN_13675 : _GEN_10603; // @[icache.scala 138:25]
  wire [184:0] _GEN_14700 = lookup & dirty ? _GEN_13676 : _GEN_10604; // @[icache.scala 138:25]
  wire [184:0] _GEN_14701 = lookup & dirty ? _GEN_13677 : _GEN_10605; // @[icache.scala 138:25]
  wire [184:0] _GEN_14702 = lookup & dirty ? _GEN_13678 : _GEN_10606; // @[icache.scala 138:25]
  wire [184:0] _GEN_14703 = lookup & dirty ? _GEN_13679 : _GEN_10607; // @[icache.scala 138:25]
  wire [184:0] _GEN_14704 = lookup & dirty ? _GEN_13680 : _GEN_10608; // @[icache.scala 138:25]
  wire [184:0] _GEN_14705 = lookup & dirty ? _GEN_13681 : _GEN_10609; // @[icache.scala 138:25]
  wire [184:0] _GEN_14706 = lookup & dirty ? _GEN_13682 : _GEN_10610; // @[icache.scala 138:25]
  wire [184:0] _GEN_14707 = lookup & dirty ? _GEN_13683 : _GEN_10611; // @[icache.scala 138:25]
  wire [184:0] _GEN_14708 = lookup & dirty ? _GEN_13684 : _GEN_10612; // @[icache.scala 138:25]
  wire [184:0] _GEN_14709 = lookup & dirty ? _GEN_13685 : _GEN_10613; // @[icache.scala 138:25]
  wire [184:0] _GEN_14710 = lookup & dirty ? _GEN_13686 : _GEN_10614; // @[icache.scala 138:25]
  wire [184:0] _GEN_14711 = lookup & dirty ? _GEN_13687 : _GEN_10615; // @[icache.scala 138:25]
  wire [184:0] _GEN_14712 = lookup & dirty ? _GEN_13688 : _GEN_10616; // @[icache.scala 138:25]
  wire [184:0] _GEN_14713 = lookup & dirty ? _GEN_13689 : _GEN_10617; // @[icache.scala 138:25]
  wire [184:0] _GEN_14714 = lookup & dirty ? _GEN_13690 : _GEN_10618; // @[icache.scala 138:25]
  wire [184:0] _GEN_14715 = lookup & dirty ? _GEN_13691 : _GEN_10619; // @[icache.scala 138:25]
  wire [184:0] _GEN_14716 = lookup & dirty ? _GEN_13692 : _GEN_10620; // @[icache.scala 138:25]
  wire [184:0] _GEN_14717 = lookup & dirty ? _GEN_13693 : _GEN_10621; // @[icache.scala 138:25]
  wire [184:0] _GEN_14718 = lookup & dirty ? _GEN_13694 : _GEN_10622; // @[icache.scala 138:25]
  wire [184:0] _GEN_14719 = lookup & dirty ? _GEN_13695 : _GEN_10623; // @[icache.scala 138:25]
  wire [184:0] _GEN_14720 = lookup & dirty ? _GEN_13696 : _GEN_10624; // @[icache.scala 138:25]
  wire [184:0] _GEN_14721 = lookup & dirty ? _GEN_13697 : _GEN_10625; // @[icache.scala 138:25]
  wire [184:0] _GEN_14722 = lookup & dirty ? _GEN_13698 : _GEN_10626; // @[icache.scala 138:25]
  wire [184:0] _GEN_14723 = lookup & dirty ? _GEN_13699 : _GEN_10627; // @[icache.scala 138:25]
  wire [184:0] _GEN_14724 = lookup & dirty ? _GEN_13700 : _GEN_10628; // @[icache.scala 138:25]
  wire [184:0] _GEN_14725 = lookup & dirty ? _GEN_13701 : _GEN_10629; // @[icache.scala 138:25]
  wire [184:0] _GEN_14726 = lookup & dirty ? _GEN_13702 : _GEN_10630; // @[icache.scala 138:25]
  wire [184:0] _GEN_14727 = lookup & dirty ? _GEN_13703 : _GEN_10631; // @[icache.scala 138:25]
  wire [184:0] _GEN_14728 = lookup & dirty ? _GEN_13704 : _GEN_10632; // @[icache.scala 138:25]
  wire [184:0] _GEN_14729 = lookup & dirty ? _GEN_13705 : _GEN_10633; // @[icache.scala 138:25]
  wire [184:0] _GEN_14730 = lookup & dirty ? _GEN_13706 : _GEN_10634; // @[icache.scala 138:25]
  wire [184:0] _GEN_14731 = lookup & dirty ? _GEN_13707 : _GEN_10635; // @[icache.scala 138:25]
  wire [184:0] _GEN_14732 = lookup & dirty ? _GEN_13708 : _GEN_10636; // @[icache.scala 138:25]
  wire [184:0] _GEN_14733 = lookup & dirty ? _GEN_13709 : _GEN_10637; // @[icache.scala 138:25]
  wire [184:0] _GEN_14734 = lookup & dirty ? _GEN_13710 : _GEN_10638; // @[icache.scala 138:25]
  wire [184:0] _GEN_14735 = lookup & dirty ? _GEN_13711 : _GEN_10639; // @[icache.scala 138:25]
  wire [184:0] _GEN_14736 = lookup & dirty ? _GEN_13712 : _GEN_10640; // @[icache.scala 138:25]
  wire [184:0] _GEN_14737 = lookup & dirty ? _GEN_13713 : _GEN_10641; // @[icache.scala 138:25]
  wire [184:0] _GEN_14738 = lookup & dirty ? _GEN_13714 : _GEN_10642; // @[icache.scala 138:25]
  wire [184:0] _GEN_14739 = lookup & dirty ? _GEN_13715 : _GEN_10643; // @[icache.scala 138:25]
  wire [184:0] _GEN_14740 = lookup & dirty ? _GEN_13716 : _GEN_10644; // @[icache.scala 138:25]
  wire [184:0] _GEN_14741 = lookup & dirty ? _GEN_13717 : _GEN_10645; // @[icache.scala 138:25]
  wire [184:0] _GEN_14742 = lookup & dirty ? _GEN_13718 : _GEN_10646; // @[icache.scala 138:25]
  wire [184:0] _GEN_14743 = lookup & dirty ? _GEN_13719 : _GEN_10647; // @[icache.scala 138:25]
  wire [184:0] _GEN_14744 = lookup & dirty ? _GEN_13720 : _GEN_10648; // @[icache.scala 138:25]
  wire [184:0] _GEN_14745 = lookup & dirty ? _GEN_13721 : _GEN_10649; // @[icache.scala 138:25]
  wire [184:0] _GEN_14746 = lookup & dirty ? _GEN_13722 : _GEN_10650; // @[icache.scala 138:25]
  wire [184:0] _GEN_14747 = lookup & dirty ? _GEN_13723 : _GEN_10651; // @[icache.scala 138:25]
  wire [184:0] _GEN_14748 = lookup & dirty ? _GEN_13724 : _GEN_10652; // @[icache.scala 138:25]
  wire [184:0] _GEN_14749 = lookup & dirty ? _GEN_13725 : _GEN_10653; // @[icache.scala 138:25]
  wire [184:0] _GEN_14750 = lookup & dirty ? _GEN_13726 : _GEN_10654; // @[icache.scala 138:25]
  wire [184:0] _GEN_14751 = lookup & dirty ? _GEN_13727 : _GEN_10655; // @[icache.scala 138:25]
  wire [184:0] _GEN_14752 = lookup & dirty ? _GEN_13728 : _GEN_10656; // @[icache.scala 138:25]
  wire [184:0] _GEN_14753 = lookup & dirty ? _GEN_13729 : _GEN_10657; // @[icache.scala 138:25]
  wire [184:0] _GEN_14754 = lookup & dirty ? _GEN_13730 : _GEN_10658; // @[icache.scala 138:25]
  wire [184:0] _GEN_14755 = lookup & dirty ? _GEN_13731 : _GEN_10659; // @[icache.scala 138:25]
  wire [184:0] _GEN_14756 = lookup & dirty ? _GEN_13732 : _GEN_10660; // @[icache.scala 138:25]
  wire [184:0] _GEN_14757 = lookup & dirty ? _GEN_13733 : _GEN_10661; // @[icache.scala 138:25]
  wire [184:0] _GEN_14758 = lookup & dirty ? _GEN_13734 : _GEN_10662; // @[icache.scala 138:25]
  wire [184:0] _GEN_14759 = lookup & dirty ? _GEN_13735 : _GEN_10663; // @[icache.scala 138:25]
  wire [184:0] _GEN_14760 = lookup & dirty ? _GEN_13736 : _GEN_10664; // @[icache.scala 138:25]
  wire [184:0] _GEN_14761 = lookup & dirty ? _GEN_13737 : _GEN_10665; // @[icache.scala 138:25]
  wire [184:0] _GEN_14762 = lookup & dirty ? _GEN_13738 : _GEN_10666; // @[icache.scala 138:25]
  wire [184:0] _GEN_14763 = lookup & dirty ? _GEN_13739 : _GEN_10667; // @[icache.scala 138:25]
  wire [184:0] _GEN_14764 = lookup & dirty ? _GEN_13740 : _GEN_10668; // @[icache.scala 138:25]
  wire [184:0] _GEN_14765 = lookup & dirty ? _GEN_13741 : _GEN_10669; // @[icache.scala 138:25]
  wire [184:0] _GEN_14766 = lookup & dirty ? _GEN_13742 : _GEN_10670; // @[icache.scala 138:25]
  wire [184:0] _GEN_14767 = lookup & dirty ? _GEN_13743 : _GEN_10671; // @[icache.scala 138:25]
  wire [184:0] _GEN_14768 = lookup & dirty ? _GEN_13744 : _GEN_10672; // @[icache.scala 138:25]
  wire [184:0] _GEN_14769 = lookup & dirty ? _GEN_13745 : _GEN_10673; // @[icache.scala 138:25]
  wire [184:0] _GEN_14770 = lookup & dirty ? _GEN_13746 : _GEN_10674; // @[icache.scala 138:25]
  wire [184:0] _GEN_14771 = lookup & dirty ? _GEN_13747 : _GEN_10675; // @[icache.scala 138:25]
  wire [184:0] _GEN_14772 = lookup & dirty ? _GEN_13748 : _GEN_10676; // @[icache.scala 138:25]
  wire [184:0] _GEN_14773 = lookup & dirty ? _GEN_13749 : _GEN_10677; // @[icache.scala 138:25]
  wire [184:0] _GEN_14774 = lookup & dirty ? _GEN_13750 : _GEN_10678; // @[icache.scala 138:25]
  wire [184:0] _GEN_14775 = lookup & dirty ? _GEN_13751 : _GEN_10679; // @[icache.scala 138:25]
  wire [184:0] _GEN_14776 = lookup & dirty ? _GEN_13752 : _GEN_10680; // @[icache.scala 138:25]
  wire [184:0] _GEN_14777 = lookup & dirty ? _GEN_13753 : _GEN_10681; // @[icache.scala 138:25]
  wire [184:0] _GEN_14778 = lookup & dirty ? _GEN_13754 : _GEN_10682; // @[icache.scala 138:25]
  wire [184:0] _GEN_14779 = lookup & dirty ? _GEN_13755 : _GEN_10683; // @[icache.scala 138:25]
  wire [184:0] _GEN_14780 = lookup & dirty ? _GEN_13756 : _GEN_10684; // @[icache.scala 138:25]
  wire [184:0] _GEN_14781 = lookup & dirty ? _GEN_13757 : _GEN_10685; // @[icache.scala 138:25]
  wire [184:0] _GEN_14782 = lookup & dirty ? _GEN_13758 : _GEN_10686; // @[icache.scala 138:25]
  wire [184:0] _GEN_14783 = lookup & dirty ? _GEN_13759 : _GEN_10687; // @[icache.scala 138:25]
  wire [184:0] _GEN_14784 = lookup & dirty ? _GEN_13760 : _GEN_10688; // @[icache.scala 138:25]
  wire [184:0] _GEN_14785 = lookup & dirty ? _GEN_13761 : _GEN_10689; // @[icache.scala 138:25]
  wire [184:0] _GEN_14786 = lookup & dirty ? _GEN_13762 : _GEN_10690; // @[icache.scala 138:25]
  wire [184:0] _GEN_14787 = lookup & dirty ? _GEN_13763 : _GEN_10691; // @[icache.scala 138:25]
  wire [184:0] _GEN_14788 = lookup & dirty ? _GEN_13764 : _GEN_10692; // @[icache.scala 138:25]
  wire [184:0] _GEN_14789 = lookup & dirty ? _GEN_13765 : _GEN_10693; // @[icache.scala 138:25]
  wire [184:0] _GEN_14790 = lookup & dirty ? _GEN_13766 : _GEN_10694; // @[icache.scala 138:25]
  wire [184:0] _GEN_14791 = lookup & dirty ? _GEN_13767 : _GEN_10695; // @[icache.scala 138:25]
  wire [184:0] _GEN_14792 = lookup & dirty ? _GEN_13768 : _GEN_10696; // @[icache.scala 138:25]
  wire [184:0] _GEN_14793 = lookup & dirty ? _GEN_13769 : _GEN_10697; // @[icache.scala 138:25]
  wire [184:0] _GEN_14794 = lookup & dirty ? _GEN_13770 : _GEN_10698; // @[icache.scala 138:25]
  wire [184:0] _GEN_14795 = lookup & dirty ? _GEN_13771 : _GEN_10699; // @[icache.scala 138:25]
  wire [184:0] _GEN_14796 = lookup & dirty ? _GEN_13772 : _GEN_10700; // @[icache.scala 138:25]
  wire [184:0] _GEN_14797 = lookup & dirty ? _GEN_13773 : _GEN_10701; // @[icache.scala 138:25]
  wire [184:0] _GEN_14798 = lookup & dirty ? _GEN_13774 : _GEN_10702; // @[icache.scala 138:25]
  wire [184:0] _GEN_14799 = lookup & dirty ? _GEN_13775 : _GEN_10703; // @[icache.scala 138:25]
  wire [184:0] _GEN_14800 = lookup & dirty ? _GEN_13776 : _GEN_10704; // @[icache.scala 138:25]
  wire [184:0] _GEN_14801 = lookup & dirty ? _GEN_13777 : _GEN_10705; // @[icache.scala 138:25]
  wire [184:0] _GEN_14802 = lookup & dirty ? _GEN_13778 : _GEN_10706; // @[icache.scala 138:25]
  wire [184:0] _GEN_14803 = lookup & dirty ? _GEN_13779 : _GEN_10707; // @[icache.scala 138:25]
  wire [184:0] _GEN_14804 = lookup & dirty ? _GEN_13780 : _GEN_10708; // @[icache.scala 138:25]
  wire [184:0] _GEN_14805 = lookup & dirty ? _GEN_13781 : _GEN_10709; // @[icache.scala 138:25]
  wire [184:0] _GEN_14806 = lookup & dirty ? _GEN_13782 : _GEN_10710; // @[icache.scala 138:25]
  wire [184:0] _GEN_14807 = lookup & dirty ? _GEN_13783 : _GEN_10711; // @[icache.scala 138:25]
  wire [184:0] _GEN_14808 = lookup & dirty ? _GEN_13784 : _GEN_10712; // @[icache.scala 138:25]
  wire [184:0] _GEN_14809 = lookup & dirty ? _GEN_13785 : _GEN_10713; // @[icache.scala 138:25]
  wire [184:0] _GEN_14810 = lookup & dirty ? _GEN_13786 : _GEN_10714; // @[icache.scala 138:25]
  wire [184:0] _GEN_14811 = lookup & dirty ? _GEN_13787 : _GEN_10715; // @[icache.scala 138:25]
  wire [184:0] _GEN_14812 = lookup & dirty ? _GEN_13788 : _GEN_10716; // @[icache.scala 138:25]
  wire [184:0] _GEN_14813 = lookup & dirty ? _GEN_13789 : _GEN_10717; // @[icache.scala 138:25]
  wire [184:0] _GEN_14814 = lookup & dirty ? _GEN_13790 : _GEN_10718; // @[icache.scala 138:25]
  wire [184:0] _GEN_14815 = lookup & dirty ? _GEN_13791 : _GEN_10719; // @[icache.scala 138:25]
  wire [184:0] _GEN_14816 = lookup & dirty ? _GEN_13792 : _GEN_10720; // @[icache.scala 138:25]
  wire [184:0] _GEN_14817 = lookup & dirty ? _GEN_13793 : _GEN_10721; // @[icache.scala 138:25]
  wire [184:0] _GEN_14818 = lookup & dirty ? _GEN_13794 : _GEN_10722; // @[icache.scala 138:25]
  wire [184:0] _GEN_14819 = lookup & dirty ? _GEN_13795 : _GEN_10723; // @[icache.scala 138:25]
  wire [184:0] _GEN_14820 = lookup & dirty ? _GEN_13796 : _GEN_10724; // @[icache.scala 138:25]
  wire [184:0] _GEN_14821 = lookup & dirty ? _GEN_13797 : _GEN_10725; // @[icache.scala 138:25]
  wire [184:0] _GEN_14822 = lookup & dirty ? _GEN_13798 : _GEN_10726; // @[icache.scala 138:25]
  wire [184:0] _GEN_14823 = lookup & dirty ? _GEN_13799 : _GEN_10727; // @[icache.scala 138:25]
  wire [184:0] _GEN_14824 = lookup & dirty ? _GEN_13800 : _GEN_10728; // @[icache.scala 138:25]
  wire [184:0] _GEN_14825 = lookup & dirty ? _GEN_13801 : _GEN_10729; // @[icache.scala 138:25]
  wire [184:0] _GEN_14826 = lookup & dirty ? _GEN_13802 : _GEN_10730; // @[icache.scala 138:25]
  wire [184:0] _GEN_14827 = lookup & dirty ? _GEN_13803 : _GEN_10731; // @[icache.scala 138:25]
  wire [184:0] _GEN_14828 = lookup & dirty ? _GEN_13804 : _GEN_10732; // @[icache.scala 138:25]
  wire [184:0] _GEN_14829 = lookup & dirty ? _GEN_13805 : _GEN_10733; // @[icache.scala 138:25]
  wire [184:0] _GEN_14830 = lookup & dirty ? _GEN_13806 : _GEN_10734; // @[icache.scala 138:25]
  wire [184:0] _GEN_14831 = lookup & dirty ? _GEN_13807 : _GEN_10735; // @[icache.scala 138:25]
  wire [184:0] _GEN_14832 = lookup & dirty ? _GEN_13808 : _GEN_10736; // @[icache.scala 138:25]
  wire [184:0] _GEN_14833 = lookup & dirty ? _GEN_13809 : _GEN_10737; // @[icache.scala 138:25]
  wire [184:0] _GEN_14834 = lookup & dirty ? _GEN_13810 : _GEN_10738; // @[icache.scala 138:25]
  wire [184:0] _GEN_14835 = lookup & dirty ? _GEN_13811 : _GEN_10739; // @[icache.scala 138:25]
  wire [184:0] _GEN_14836 = lookup & dirty ? _GEN_13812 : _GEN_10740; // @[icache.scala 138:25]
  wire [184:0] _GEN_14837 = lookup & dirty ? _GEN_13813 : _GEN_10741; // @[icache.scala 138:25]
  wire [184:0] _GEN_14838 = lookup & dirty ? _GEN_13814 : _GEN_10742; // @[icache.scala 138:25]
  wire [184:0] _GEN_14839 = lookup & dirty ? _GEN_13815 : _GEN_10743; // @[icache.scala 138:25]
  wire [184:0] _GEN_14840 = lookup & dirty ? _GEN_13816 : _GEN_10744; // @[icache.scala 138:25]
  wire [184:0] _GEN_14841 = lookup & dirty ? _GEN_13817 : _GEN_10745; // @[icache.scala 138:25]
  wire [184:0] _GEN_14842 = lookup & dirty ? _GEN_13818 : _GEN_10746; // @[icache.scala 138:25]
  wire [184:0] _GEN_14843 = lookup & dirty ? _GEN_13819 : _GEN_10747; // @[icache.scala 138:25]
  wire [184:0] _GEN_14844 = lookup & dirty ? _GEN_13820 : _GEN_10748; // @[icache.scala 138:25]
  wire [184:0] _GEN_14845 = lookup & dirty ? _GEN_13821 : _GEN_10749; // @[icache.scala 138:25]
  wire [184:0] _GEN_14846 = lookup & dirty ? _GEN_13822 : _GEN_10750; // @[icache.scala 138:25]
  wire [184:0] _GEN_14847 = lookup & dirty ? _GEN_13823 : _GEN_10751; // @[icache.scala 138:25]
  wire [184:0] _GEN_14848 = lookup & dirty ? _GEN_13824 : _GEN_10752; // @[icache.scala 138:25]
  wire [184:0] _GEN_14849 = lookup & dirty ? _GEN_13825 : _GEN_10753; // @[icache.scala 138:25]
  wire [184:0] _GEN_14850 = lookup & dirty ? _GEN_13826 : _GEN_10754; // @[icache.scala 138:25]
  wire [184:0] _GEN_14851 = lookup & dirty ? _GEN_13827 : _GEN_10755; // @[icache.scala 138:25]
  wire [184:0] _GEN_14852 = lookup & dirty ? _GEN_13828 : _GEN_10756; // @[icache.scala 138:25]
  wire [184:0] _GEN_14853 = lookup & dirty ? _GEN_13829 : _GEN_10757; // @[icache.scala 138:25]
  wire [184:0] _GEN_14854 = lookup & dirty ? _GEN_13830 : _GEN_10758; // @[icache.scala 138:25]
  wire [184:0] _GEN_14855 = lookup & dirty ? _GEN_13831 : _GEN_10759; // @[icache.scala 138:25]
  wire [184:0] _GEN_14856 = lookup & dirty ? _GEN_13832 : _GEN_10760; // @[icache.scala 138:25]
  wire [184:0] _GEN_14857 = lookup & dirty ? _GEN_13833 : _GEN_10761; // @[icache.scala 138:25]
  wire [184:0] _GEN_14858 = lookup & dirty ? _GEN_13834 : _GEN_10762; // @[icache.scala 138:25]
  wire [184:0] _GEN_14859 = lookup & dirty ? _GEN_13835 : _GEN_10763; // @[icache.scala 138:25]
  wire [184:0] _GEN_14860 = lookup & dirty ? _GEN_13836 : _GEN_10764; // @[icache.scala 138:25]
  wire [184:0] _GEN_14861 = lookup & dirty ? _GEN_13837 : _GEN_10765; // @[icache.scala 138:25]
  wire [184:0] _GEN_14862 = lookup & dirty ? _GEN_13838 : _GEN_10766; // @[icache.scala 138:25]
  wire [184:0] _GEN_14863 = lookup & dirty ? _GEN_13839 : _GEN_10767; // @[icache.scala 138:25]
  wire [184:0] _GEN_14864 = lookup & dirty ? _GEN_13840 : _GEN_10768; // @[icache.scala 138:25]
  wire [184:0] _GEN_14865 = lookup & dirty ? _GEN_13841 : _GEN_10769; // @[icache.scala 138:25]
  wire [184:0] _GEN_14866 = lookup & dirty ? _GEN_13842 : _GEN_10770; // @[icache.scala 138:25]
  wire [184:0] _GEN_14867 = lookup & dirty ? _GEN_13843 : _GEN_10771; // @[icache.scala 138:25]
  wire [184:0] _GEN_14868 = lookup & dirty ? _GEN_13844 : _GEN_10772; // @[icache.scala 138:25]
  wire [184:0] _GEN_14869 = lookup & dirty ? _GEN_13845 : _GEN_10773; // @[icache.scala 138:25]
  wire [184:0] _GEN_14870 = lookup & dirty ? _GEN_13846 : _GEN_10774; // @[icache.scala 138:25]
  wire [184:0] _GEN_14871 = lookup & dirty ? _GEN_13847 : _GEN_10775; // @[icache.scala 138:25]
  wire [184:0] _GEN_14872 = lookup & dirty ? _GEN_13848 : _GEN_10776; // @[icache.scala 138:25]
  wire [184:0] _GEN_14873 = lookup & dirty ? _GEN_13849 : _GEN_10777; // @[icache.scala 138:25]
  wire [184:0] _GEN_14874 = lookup & dirty ? _GEN_13850 : _GEN_10778; // @[icache.scala 138:25]
  wire [184:0] _GEN_14875 = lookup & dirty ? _GEN_13851 : _GEN_10779; // @[icache.scala 138:25]
  wire [184:0] _GEN_14876 = lookup & dirty ? _GEN_13852 : _GEN_10780; // @[icache.scala 138:25]
  wire [184:0] _GEN_14877 = lookup & dirty ? _GEN_13853 : _GEN_10781; // @[icache.scala 138:25]
  wire [184:0] _GEN_14878 = lookup & dirty ? _GEN_13854 : _GEN_10782; // @[icache.scala 138:25]
  wire [184:0] _GEN_14879 = lookup & dirty ? _GEN_13855 : _GEN_10783; // @[icache.scala 138:25]
  wire [184:0] _GEN_14880 = lookup & dirty ? _GEN_13856 : _GEN_10784; // @[icache.scala 138:25]
  wire [184:0] _GEN_14881 = lookup & dirty ? _GEN_13857 : _GEN_10785; // @[icache.scala 138:25]
  wire [184:0] _GEN_14882 = lookup & dirty ? _GEN_13858 : _GEN_10786; // @[icache.scala 138:25]
  wire [184:0] _GEN_14883 = lookup & dirty ? _GEN_13859 : _GEN_10787; // @[icache.scala 138:25]
  wire [184:0] _GEN_14884 = lookup & dirty ? _GEN_13860 : _GEN_10788; // @[icache.scala 138:25]
  wire [184:0] _GEN_14885 = lookup & dirty ? _GEN_13861 : _GEN_10789; // @[icache.scala 138:25]
  wire [184:0] _GEN_14886 = lookup & dirty ? _GEN_13862 : _GEN_10790; // @[icache.scala 138:25]
  wire [184:0] _GEN_14887 = lookup & dirty ? _GEN_13863 : _GEN_10791; // @[icache.scala 138:25]
  wire [184:0] _GEN_14888 = lookup & dirty ? _GEN_13864 : _GEN_10792; // @[icache.scala 138:25]
  wire [184:0] _GEN_14889 = lookup & dirty ? _GEN_13865 : _GEN_10793; // @[icache.scala 138:25]
  wire [184:0] _GEN_14890 = lookup & dirty ? _GEN_13866 : _GEN_10794; // @[icache.scala 138:25]
  wire [184:0] _GEN_14891 = lookup & dirty ? _GEN_13867 : _GEN_10795; // @[icache.scala 138:25]
  wire [184:0] _GEN_14892 = lookup & dirty ? _GEN_13868 : _GEN_10796; // @[icache.scala 138:25]
  wire [184:0] _GEN_14893 = lookup & dirty ? _GEN_13869 : _GEN_10797; // @[icache.scala 138:25]
  wire [184:0] _GEN_14894 = lookup & dirty ? _GEN_13870 : _GEN_10798; // @[icache.scala 138:25]
  wire [184:0] _GEN_14895 = lookup & dirty ? _GEN_13871 : _GEN_10799; // @[icache.scala 138:25]
  wire [184:0] _GEN_14896 = lookup & dirty ? _GEN_13872 : _GEN_10800; // @[icache.scala 138:25]
  wire [184:0] _GEN_14897 = lookup & dirty ? _GEN_13873 : _GEN_10801; // @[icache.scala 138:25]
  wire [184:0] _GEN_14898 = lookup & dirty ? _GEN_13874 : _GEN_10802; // @[icache.scala 138:25]
  wire [184:0] _GEN_14899 = lookup & dirty ? _GEN_13875 : _GEN_10803; // @[icache.scala 138:25]
  wire [184:0] _GEN_14900 = lookup & dirty ? _GEN_13876 : _GEN_10804; // @[icache.scala 138:25]
  wire [184:0] _GEN_14901 = lookup & dirty ? _GEN_13877 : _GEN_10805; // @[icache.scala 138:25]
  wire [184:0] _GEN_14902 = lookup & dirty ? _GEN_13878 : _GEN_10806; // @[icache.scala 138:25]
  wire [184:0] _GEN_14903 = lookup & dirty ? _GEN_13879 : _GEN_10807; // @[icache.scala 138:25]
  wire [184:0] _GEN_14904 = lookup & dirty ? _GEN_13880 : _GEN_10808; // @[icache.scala 138:25]
  wire [184:0] _GEN_14905 = lookup & dirty ? _GEN_13881 : _GEN_10809; // @[icache.scala 138:25]
  wire [184:0] _GEN_14906 = lookup & dirty ? _GEN_13882 : _GEN_10810; // @[icache.scala 138:25]
  wire [184:0] _GEN_14907 = lookup & dirty ? _GEN_13883 : _GEN_10811; // @[icache.scala 138:25]
  wire [184:0] _GEN_14908 = lookup & dirty ? _GEN_13884 : _GEN_10812; // @[icache.scala 138:25]
  wire [184:0] _GEN_14909 = lookup & dirty ? _GEN_13885 : _GEN_10813; // @[icache.scala 138:25]
  wire [184:0] _GEN_14910 = lookup & dirty ? _GEN_13886 : _GEN_10814; // @[icache.scala 138:25]
  wire [184:0] _GEN_14911 = lookup & dirty ? _GEN_13887 : _GEN_10815; // @[icache.scala 138:25]
  wire [184:0] _GEN_14912 = lookup & dirty ? _GEN_13888 : _GEN_10816; // @[icache.scala 138:25]
  wire [184:0] _GEN_14913 = lookup & dirty ? _GEN_13889 : _GEN_10817; // @[icache.scala 138:25]
  wire [184:0] _GEN_14914 = lookup & dirty ? _GEN_13890 : _GEN_10818; // @[icache.scala 138:25]
  wire [184:0] _GEN_14915 = lookup & dirty ? _GEN_13891 : _GEN_10819; // @[icache.scala 138:25]
  wire [184:0] _GEN_14916 = lookup & dirty ? _GEN_13892 : _GEN_10820; // @[icache.scala 138:25]
  wire [184:0] _GEN_14917 = lookup & dirty ? _GEN_13893 : _GEN_10821; // @[icache.scala 138:25]
  wire [184:0] _GEN_14918 = lookup & dirty ? _GEN_13894 : _GEN_10822; // @[icache.scala 138:25]
  wire [184:0] _GEN_14919 = lookup & dirty ? _GEN_13895 : _GEN_10823; // @[icache.scala 138:25]
  wire [184:0] _GEN_14920 = lookup & dirty ? _GEN_13896 : _GEN_10824; // @[icache.scala 138:25]
  wire [184:0] _GEN_14921 = lookup & dirty ? _GEN_13897 : _GEN_10825; // @[icache.scala 138:25]
  wire [184:0] _GEN_14922 = lookup & dirty ? _GEN_13898 : _GEN_10826; // @[icache.scala 138:25]
  wire [184:0] _GEN_14923 = lookup & dirty ? _GEN_13899 : _GEN_10827; // @[icache.scala 138:25]
  wire [184:0] _GEN_14924 = lookup & dirty ? _GEN_13900 : _GEN_10828; // @[icache.scala 138:25]
  wire [184:0] _GEN_14925 = lookup & dirty ? _GEN_13901 : _GEN_10829; // @[icache.scala 138:25]
  wire [184:0] _GEN_14926 = lookup & dirty ? _GEN_13902 : _GEN_10830; // @[icache.scala 138:25]
  wire [184:0] _GEN_14927 = lookup & dirty ? _GEN_13903 : _GEN_10831; // @[icache.scala 138:25]
  wire [184:0] _GEN_14928 = lookup & dirty ? _GEN_13904 : _GEN_10832; // @[icache.scala 138:25]
  wire [184:0] _GEN_14929 = lookup & dirty ? _GEN_13905 : _GEN_10833; // @[icache.scala 138:25]
  wire [184:0] _GEN_14930 = lookup & dirty ? _GEN_13906 : _GEN_10834; // @[icache.scala 138:25]
  wire [184:0] _GEN_14931 = lookup & dirty ? _GEN_13907 : _GEN_10835; // @[icache.scala 138:25]
  wire [184:0] _GEN_14932 = lookup & dirty ? _GEN_13908 : _GEN_10836; // @[icache.scala 138:25]
  wire [184:0] _GEN_14933 = lookup & dirty ? _GEN_13909 : _GEN_10837; // @[icache.scala 138:25]
  wire [184:0] _GEN_14934 = lookup & dirty ? _GEN_13910 : _GEN_10838; // @[icache.scala 138:25]
  wire [184:0] _GEN_14935 = lookup & dirty ? _GEN_13911 : _GEN_10839; // @[icache.scala 138:25]
  wire [184:0] _GEN_14936 = lookup & dirty ? _GEN_13912 : _GEN_10840; // @[icache.scala 138:25]
  wire [184:0] _GEN_14937 = lookup & dirty ? _GEN_13913 : _GEN_10841; // @[icache.scala 138:25]
  wire [184:0] _GEN_14938 = lookup & dirty ? _GEN_13914 : _GEN_10842; // @[icache.scala 138:25]
  wire [184:0] _GEN_14939 = lookup & dirty ? _GEN_13915 : _GEN_10843; // @[icache.scala 138:25]
  wire [184:0] _GEN_14940 = lookup & dirty ? _GEN_13916 : _GEN_10844; // @[icache.scala 138:25]
  wire [184:0] _GEN_14941 = lookup & dirty ? _GEN_13917 : _GEN_10845; // @[icache.scala 138:25]
  wire [184:0] _GEN_14942 = lookup & dirty ? _GEN_13918 : _GEN_10846; // @[icache.scala 138:25]
  wire [184:0] _GEN_14943 = lookup & dirty ? _GEN_13919 : _GEN_10847; // @[icache.scala 138:25]
  wire [184:0] _GEN_14944 = lookup & dirty ? _GEN_13920 : _GEN_10848; // @[icache.scala 138:25]
  wire [184:0] _GEN_14945 = lookup & dirty ? _GEN_13921 : _GEN_10849; // @[icache.scala 138:25]
  wire [184:0] _GEN_14946 = lookup & dirty ? _GEN_13922 : _GEN_10850; // @[icache.scala 138:25]
  wire [184:0] _GEN_14947 = lookup & dirty ? _GEN_13923 : _GEN_10851; // @[icache.scala 138:25]
  wire [184:0] _GEN_14948 = lookup & dirty ? _GEN_13924 : _GEN_10852; // @[icache.scala 138:25]
  wire [184:0] _GEN_14949 = lookup & dirty ? _GEN_13925 : _GEN_10853; // @[icache.scala 138:25]
  wire [184:0] _GEN_14950 = lookup & dirty ? _GEN_13926 : _GEN_10854; // @[icache.scala 138:25]
  wire [184:0] _GEN_14951 = lookup & dirty ? _GEN_13927 : _GEN_10855; // @[icache.scala 138:25]
  wire [184:0] _GEN_14952 = lookup & dirty ? _GEN_13928 : _GEN_10856; // @[icache.scala 138:25]
  wire [184:0] _GEN_14953 = lookup & dirty ? _GEN_13929 : _GEN_10857; // @[icache.scala 138:25]
  wire [184:0] _GEN_14954 = lookup & dirty ? _GEN_13930 : _GEN_10858; // @[icache.scala 138:25]
  wire [184:0] _GEN_14955 = lookup & dirty ? _GEN_13931 : _GEN_10859; // @[icache.scala 138:25]
  wire [184:0] _GEN_14956 = lookup & dirty ? _GEN_13932 : _GEN_10860; // @[icache.scala 138:25]
  wire [184:0] _GEN_14957 = lookup & dirty ? _GEN_13933 : _GEN_10861; // @[icache.scala 138:25]
  wire [184:0] _GEN_14958 = lookup & dirty ? _GEN_13934 : _GEN_10862; // @[icache.scala 138:25]
  wire [184:0] _GEN_14959 = lookup & dirty ? _GEN_13935 : _GEN_10863; // @[icache.scala 138:25]
  wire [184:0] _GEN_14960 = lookup & dirty ? _GEN_13936 : _GEN_10864; // @[icache.scala 138:25]
  wire [184:0] _GEN_14961 = lookup & dirty ? _GEN_13937 : _GEN_10865; // @[icache.scala 138:25]
  wire [184:0] _GEN_14962 = lookup & dirty ? _GEN_13938 : _GEN_10866; // @[icache.scala 138:25]
  wire [184:0] _GEN_14963 = lookup & dirty ? _GEN_13939 : _GEN_10867; // @[icache.scala 138:25]
  wire [184:0] _GEN_14964 = lookup & dirty ? _GEN_13940 : _GEN_10868; // @[icache.scala 138:25]
  wire [184:0] _GEN_14965 = lookup & dirty ? _GEN_13941 : _GEN_10869; // @[icache.scala 138:25]
  wire [184:0] _GEN_14966 = lookup & dirty ? _GEN_13942 : _GEN_10870; // @[icache.scala 138:25]
  wire [184:0] _GEN_14967 = lookup & dirty ? _GEN_13943 : _GEN_10871; // @[icache.scala 138:25]
  wire [184:0] _GEN_14968 = lookup & dirty ? _GEN_13944 : _GEN_10872; // @[icache.scala 138:25]
  wire [184:0] _GEN_14969 = lookup & dirty ? _GEN_13945 : _GEN_10873; // @[icache.scala 138:25]
  wire [184:0] _GEN_14970 = lookup & dirty ? _GEN_13946 : _GEN_10874; // @[icache.scala 138:25]
  wire [184:0] _GEN_14971 = lookup & dirty ? _GEN_13947 : _GEN_10875; // @[icache.scala 138:25]
  wire [184:0] _GEN_14972 = lookup & dirty ? _GEN_13948 : _GEN_10876; // @[icache.scala 138:25]
  wire [184:0] _GEN_14973 = lookup & dirty ? _GEN_13949 : _GEN_10877; // @[icache.scala 138:25]
  wire [184:0] _GEN_14974 = lookup & dirty ? _GEN_13950 : _GEN_10878; // @[icache.scala 138:25]
  wire [184:0] _GEN_14975 = lookup & dirty ? _GEN_13951 : _GEN_10879; // @[icache.scala 138:25]
  wire [184:0] _GEN_14976 = lookup & dirty ? _GEN_13952 : _GEN_10880; // @[icache.scala 138:25]
  wire [184:0] _GEN_14977 = lookup & dirty ? _GEN_13953 : _GEN_10881; // @[icache.scala 138:25]
  wire [184:0] _GEN_14978 = lookup & dirty ? _GEN_13954 : _GEN_10882; // @[icache.scala 138:25]
  wire [184:0] _GEN_14979 = lookup & dirty ? _GEN_13955 : _GEN_10883; // @[icache.scala 138:25]
  wire [184:0] _GEN_14980 = lookup & dirty ? _GEN_13956 : _GEN_10884; // @[icache.scala 138:25]
  wire [184:0] _GEN_14981 = lookup & dirty ? _GEN_13957 : _GEN_10885; // @[icache.scala 138:25]
  wire [184:0] _GEN_14982 = lookup & dirty ? _GEN_13958 : _GEN_10886; // @[icache.scala 138:25]
  wire [184:0] _GEN_14983 = lookup & dirty ? _GEN_13959 : _GEN_10887; // @[icache.scala 138:25]
  wire [184:0] _GEN_14984 = lookup & dirty ? _GEN_13960 : _GEN_10888; // @[icache.scala 138:25]
  wire [184:0] _GEN_14985 = lookup & dirty ? _GEN_13961 : _GEN_10889; // @[icache.scala 138:25]
  wire [184:0] _GEN_14986 = lookup & dirty ? _GEN_13962 : _GEN_10890; // @[icache.scala 138:25]
  wire [184:0] _GEN_14987 = lookup & dirty ? _GEN_13963 : _GEN_10891; // @[icache.scala 138:25]
  wire [184:0] _GEN_14988 = lookup & dirty ? _GEN_13964 : _GEN_10892; // @[icache.scala 138:25]
  wire [184:0] _GEN_14989 = lookup & dirty ? _GEN_13965 : _GEN_10893; // @[icache.scala 138:25]
  wire [184:0] _GEN_14990 = lookup & dirty ? _GEN_13966 : _GEN_10894; // @[icache.scala 138:25]
  wire [184:0] _GEN_14991 = lookup & dirty ? _GEN_13967 : _GEN_10895; // @[icache.scala 138:25]
  wire [184:0] _GEN_14992 = lookup & dirty ? _GEN_13968 : _GEN_10896; // @[icache.scala 138:25]
  wire [184:0] _GEN_14993 = lookup & dirty ? _GEN_13969 : _GEN_10897; // @[icache.scala 138:25]
  wire [184:0] _GEN_14994 = lookup & dirty ? _GEN_13970 : _GEN_10898; // @[icache.scala 138:25]
  wire [184:0] _GEN_14995 = lookup & dirty ? _GEN_13971 : _GEN_10899; // @[icache.scala 138:25]
  wire [184:0] _GEN_14996 = lookup & dirty ? _GEN_13972 : _GEN_10900; // @[icache.scala 138:25]
  wire [184:0] _GEN_14997 = lookup & dirty ? _GEN_13973 : _GEN_10901; // @[icache.scala 138:25]
  wire [184:0] _GEN_14998 = lookup & dirty ? _GEN_13974 : _GEN_10902; // @[icache.scala 138:25]
  wire [184:0] _GEN_14999 = lookup & dirty ? _GEN_13975 : _GEN_10903; // @[icache.scala 138:25]
  wire [184:0] _GEN_15000 = lookup & dirty ? _GEN_13976 : _GEN_10904; // @[icache.scala 138:25]
  wire [184:0] _GEN_15001 = lookup & dirty ? _GEN_13977 : _GEN_10905; // @[icache.scala 138:25]
  wire [184:0] _GEN_15002 = lookup & dirty ? _GEN_13978 : _GEN_10906; // @[icache.scala 138:25]
  wire [184:0] _GEN_15003 = lookup & dirty ? _GEN_13979 : _GEN_10907; // @[icache.scala 138:25]
  wire [184:0] _GEN_15004 = lookup & dirty ? _GEN_13980 : _GEN_10908; // @[icache.scala 138:25]
  wire [184:0] _GEN_15005 = lookup & dirty ? _GEN_13981 : _GEN_10909; // @[icache.scala 138:25]
  wire [184:0] _GEN_15006 = lookup & dirty ? _GEN_13982 : _GEN_10910; // @[icache.scala 138:25]
  wire [184:0] _GEN_15007 = lookup & dirty ? _GEN_13983 : _GEN_10911; // @[icache.scala 138:25]
  wire [184:0] _GEN_15008 = lookup & dirty ? _GEN_13984 : _GEN_10912; // @[icache.scala 138:25]
  wire [184:0] _GEN_15009 = lookup & dirty ? _GEN_13985 : _GEN_10913; // @[icache.scala 138:25]
  wire [184:0] _GEN_15010 = lookup & dirty ? _GEN_13986 : _GEN_10914; // @[icache.scala 138:25]
  wire [184:0] _GEN_15011 = lookup & dirty ? _GEN_13987 : _GEN_10915; // @[icache.scala 138:25]
  wire [184:0] _GEN_15012 = lookup & dirty ? _GEN_13988 : _GEN_10916; // @[icache.scala 138:25]
  wire [184:0] _GEN_15013 = lookup & dirty ? _GEN_13989 : _GEN_10917; // @[icache.scala 138:25]
  wire [184:0] _GEN_15014 = lookup & dirty ? _GEN_13990 : _GEN_10918; // @[icache.scala 138:25]
  wire [184:0] _GEN_15015 = lookup & dirty ? _GEN_13991 : _GEN_10919; // @[icache.scala 138:25]
  wire [184:0] _GEN_15016 = lookup & dirty ? _GEN_13992 : _GEN_10920; // @[icache.scala 138:25]
  wire [184:0] _GEN_15017 = lookup & dirty ? _GEN_13993 : _GEN_10921; // @[icache.scala 138:25]
  wire [184:0] _GEN_15018 = lookup & dirty ? _GEN_13994 : _GEN_10922; // @[icache.scala 138:25]
  wire [184:0] _GEN_15019 = lookup & dirty ? _GEN_13995 : _GEN_10923; // @[icache.scala 138:25]
  wire [184:0] _GEN_15020 = lookup & dirty ? _GEN_13996 : _GEN_10924; // @[icache.scala 138:25]
  wire [184:0] _GEN_15021 = lookup & dirty ? _GEN_13997 : _GEN_10925; // @[icache.scala 138:25]
  wire [184:0] _GEN_15022 = lookup & dirty ? _GEN_13998 : _GEN_10926; // @[icache.scala 138:25]
  wire [184:0] _GEN_15023 = lookup & dirty ? _GEN_13999 : _GEN_10927; // @[icache.scala 138:25]
  wire [184:0] _GEN_15024 = lookup & dirty ? _GEN_14000 : _GEN_10928; // @[icache.scala 138:25]
  wire [184:0] _GEN_15025 = lookup & dirty ? _GEN_14001 : _GEN_10929; // @[icache.scala 138:25]
  wire [184:0] _GEN_15026 = lookup & dirty ? _GEN_14002 : _GEN_10930; // @[icache.scala 138:25]
  wire [184:0] _GEN_15027 = lookup & dirty ? _GEN_14003 : _GEN_10931; // @[icache.scala 138:25]
  wire [184:0] _GEN_15028 = lookup & dirty ? _GEN_14004 : _GEN_10932; // @[icache.scala 138:25]
  wire [184:0] _GEN_15029 = lookup & dirty ? _GEN_14005 : _GEN_10933; // @[icache.scala 138:25]
  wire [184:0] _GEN_15030 = lookup & dirty ? _GEN_14006 : _GEN_10934; // @[icache.scala 138:25]
  wire [184:0] _GEN_15031 = lookup & dirty ? _GEN_14007 : _GEN_10935; // @[icache.scala 138:25]
  wire [184:0] _GEN_15032 = lookup & dirty ? _GEN_14008 : _GEN_10936; // @[icache.scala 138:25]
  wire [184:0] _GEN_15033 = lookup & dirty ? _GEN_14009 : _GEN_10937; // @[icache.scala 138:25]
  wire [184:0] _GEN_15034 = lookup & dirty ? _GEN_14010 : _GEN_10938; // @[icache.scala 138:25]
  wire [184:0] _GEN_15035 = lookup & dirty ? _GEN_14011 : _GEN_10939; // @[icache.scala 138:25]
  wire [184:0] _GEN_15036 = lookup & dirty ? _GEN_14012 : _GEN_10940; // @[icache.scala 138:25]
  wire [184:0] _GEN_15037 = lookup & dirty ? _GEN_14013 : _GEN_10941; // @[icache.scala 138:25]
  wire [184:0] _GEN_15038 = lookup & dirty ? _GEN_14014 : _GEN_10942; // @[icache.scala 138:25]
  wire [184:0] _GEN_15039 = lookup & dirty ? _GEN_14015 : _GEN_10943; // @[icache.scala 138:25]
  wire [184:0] _GEN_15040 = lookup & dirty ? _GEN_14016 : _GEN_10944; // @[icache.scala 138:25]
  wire [184:0] _GEN_15041 = lookup & dirty ? _GEN_14017 : _GEN_10945; // @[icache.scala 138:25]
  wire [184:0] _GEN_15042 = lookup & dirty ? _GEN_14018 : _GEN_10946; // @[icache.scala 138:25]
  wire [184:0] _GEN_15043 = lookup & dirty ? _GEN_14019 : _GEN_10947; // @[icache.scala 138:25]
  wire [184:0] _GEN_15044 = lookup & dirty ? _GEN_14020 : _GEN_10948; // @[icache.scala 138:25]
  wire [184:0] _GEN_15045 = lookup & dirty ? _GEN_14021 : _GEN_10949; // @[icache.scala 138:25]
  wire [184:0] _GEN_15046 = lookup & dirty ? _GEN_14022 : _GEN_10950; // @[icache.scala 138:25]
  wire [184:0] _GEN_15047 = lookup & dirty ? _GEN_14023 : _GEN_10951; // @[icache.scala 138:25]
  wire [184:0] _GEN_15048 = lookup & dirty ? _GEN_14024 : _GEN_10952; // @[icache.scala 138:25]
  wire [184:0] _GEN_15049 = lookup & dirty ? _GEN_14025 : _GEN_10953; // @[icache.scala 138:25]
  wire [184:0] _GEN_15050 = lookup & dirty ? _GEN_14026 : _GEN_10954; // @[icache.scala 138:25]
  wire [184:0] _GEN_15051 = lookup & dirty ? _GEN_14027 : _GEN_10955; // @[icache.scala 138:25]
  wire [184:0] _GEN_15052 = lookup & dirty ? _GEN_14028 : _GEN_10956; // @[icache.scala 138:25]
  wire [184:0] _GEN_15053 = lookup & dirty ? _GEN_14029 : _GEN_10957; // @[icache.scala 138:25]
  wire [184:0] _GEN_15054 = lookup & dirty ? _GEN_14030 : _GEN_10958; // @[icache.scala 138:25]
  wire [184:0] _GEN_15055 = lookup & dirty ? _GEN_14031 : _GEN_10959; // @[icache.scala 138:25]
  wire [184:0] _GEN_15056 = lookup & dirty ? _GEN_14032 : _GEN_10960; // @[icache.scala 138:25]
  wire [184:0] _GEN_15057 = lookup & dirty ? _GEN_14033 : _GEN_10961; // @[icache.scala 138:25]
  wire [184:0] _GEN_15058 = lookup & dirty ? _GEN_14034 : _GEN_10962; // @[icache.scala 138:25]
  wire [184:0] _GEN_15059 = lookup & dirty ? _GEN_14035 : _GEN_10963; // @[icache.scala 138:25]
  wire [184:0] _GEN_15060 = lookup & dirty ? _GEN_14036 : _GEN_10964; // @[icache.scala 138:25]
  wire [184:0] _GEN_15061 = lookup & dirty ? _GEN_14037 : _GEN_10965; // @[icache.scala 138:25]
  wire [184:0] _GEN_15062 = lookup & dirty ? _GEN_14038 : _GEN_10966; // @[icache.scala 138:25]
  wire [184:0] _GEN_15063 = lookup & dirty ? _GEN_14039 : _GEN_10967; // @[icache.scala 138:25]
  wire [184:0] _GEN_15064 = lookup & dirty ? _GEN_14040 : _GEN_10968; // @[icache.scala 138:25]
  wire [184:0] _GEN_15065 = lookup & dirty ? _GEN_14041 : _GEN_10969; // @[icache.scala 138:25]
  wire [184:0] _GEN_15066 = lookup & dirty ? _GEN_14042 : _GEN_10970; // @[icache.scala 138:25]
  wire [184:0] _GEN_15067 = lookup & dirty ? _GEN_14043 : _GEN_10971; // @[icache.scala 138:25]
  wire [184:0] _GEN_15068 = lookup & dirty ? _GEN_14044 : _GEN_10972; // @[icache.scala 138:25]
  wire [184:0] _GEN_15069 = lookup & dirty ? _GEN_14045 : _GEN_10973; // @[icache.scala 138:25]
  wire [184:0] _GEN_15070 = lookup & dirty ? _GEN_14046 : _GEN_10974; // @[icache.scala 138:25]
  wire [184:0] _GEN_15071 = lookup & dirty ? _GEN_14047 : _GEN_10975; // @[icache.scala 138:25]
  wire [184:0] _GEN_15072 = lookup & dirty ? _GEN_14048 : _GEN_10976; // @[icache.scala 138:25]
  wire [184:0] _GEN_15073 = lookup & dirty ? _GEN_14049 : _GEN_10977; // @[icache.scala 138:25]
  wire [184:0] _GEN_15074 = lookup & dirty ? _GEN_14050 : _GEN_10978; // @[icache.scala 138:25]
  wire [184:0] _GEN_15075 = lookup & dirty ? _GEN_14051 : _GEN_10979; // @[icache.scala 138:25]
  wire [184:0] _GEN_15076 = lookup & dirty ? _GEN_14052 : _GEN_10980; // @[icache.scala 138:25]
  wire [184:0] _GEN_15077 = lookup & dirty ? _GEN_14053 : _GEN_10981; // @[icache.scala 138:25]
  wire [184:0] _GEN_15078 = lookup & dirty ? _GEN_14054 : _GEN_10982; // @[icache.scala 138:25]
  wire [184:0] _GEN_15079 = lookup & dirty ? _GEN_14055 : _GEN_10983; // @[icache.scala 138:25]
  wire [184:0] _GEN_15080 = lookup & dirty ? _GEN_14056 : _GEN_10984; // @[icache.scala 138:25]
  wire [184:0] _GEN_15081 = lookup & dirty ? _GEN_14057 : _GEN_10985; // @[icache.scala 138:25]
  wire [184:0] _GEN_15082 = lookup & dirty ? _GEN_14058 : _GEN_10986; // @[icache.scala 138:25]
  wire [184:0] _GEN_15083 = lookup & dirty ? _GEN_14059 : _GEN_10987; // @[icache.scala 138:25]
  wire [184:0] _GEN_15084 = lookup & dirty ? _GEN_14060 : _GEN_10988; // @[icache.scala 138:25]
  wire [184:0] _GEN_15085 = lookup & dirty ? _GEN_14061 : _GEN_10989; // @[icache.scala 138:25]
  wire [184:0] _GEN_15086 = lookup & dirty ? _GEN_14062 : _GEN_10990; // @[icache.scala 138:25]
  wire [184:0] _GEN_15087 = lookup & dirty ? _GEN_14063 : _GEN_10991; // @[icache.scala 138:25]
  wire [184:0] _GEN_15088 = lookup & dirty ? _GEN_14064 : _GEN_10992; // @[icache.scala 138:25]
  wire [184:0] _GEN_15089 = lookup & dirty ? _GEN_14065 : _GEN_10993; // @[icache.scala 138:25]
  wire [184:0] _GEN_15090 = lookup & dirty ? _GEN_14066 : _GEN_10994; // @[icache.scala 138:25]
  wire [184:0] _GEN_15091 = lookup & dirty ? _GEN_14067 : _GEN_10995; // @[icache.scala 138:25]
  wire [184:0] _GEN_15092 = lookup & dirty ? _GEN_14068 : _GEN_10996; // @[icache.scala 138:25]
  wire [184:0] _GEN_15093 = lookup & dirty ? _GEN_14069 : _GEN_10997; // @[icache.scala 138:25]
  wire [184:0] _GEN_15094 = lookup & dirty ? _GEN_14070 : _GEN_10998; // @[icache.scala 138:25]
  wire [184:0] _GEN_15095 = lookup & dirty ? _GEN_14071 : _GEN_10999; // @[icache.scala 138:25]
  wire [184:0] _GEN_15096 = lookup & dirty ? _GEN_14072 : _GEN_11000; // @[icache.scala 138:25]
  wire [184:0] _GEN_15097 = lookup & dirty ? _GEN_14073 : _GEN_11001; // @[icache.scala 138:25]
  wire [184:0] _GEN_15098 = lookup & dirty ? _GEN_14074 : _GEN_11002; // @[icache.scala 138:25]
  wire [184:0] _GEN_15099 = lookup & dirty ? _GEN_14075 : _GEN_11003; // @[icache.scala 138:25]
  wire [184:0] _GEN_15100 = lookup & dirty ? _GEN_14076 : _GEN_11004; // @[icache.scala 138:25]
  wire [184:0] _GEN_15101 = lookup & dirty ? _GEN_14077 : _GEN_11005; // @[icache.scala 138:25]
  wire [184:0] _GEN_15102 = lookup & dirty ? _GEN_14078 : _GEN_11006; // @[icache.scala 138:25]
  wire [184:0] _GEN_15103 = lookup & dirty ? _GEN_14079 : _GEN_11007; // @[icache.scala 138:25]
  wire [184:0] _GEN_15104 = lookup & dirty ? _GEN_14080 : _GEN_11008; // @[icache.scala 138:25]
  wire [184:0] _GEN_15105 = lookup & dirty ? _GEN_14081 : _GEN_11009; // @[icache.scala 138:25]
  wire [184:0] _GEN_15106 = lookup & dirty ? _GEN_14082 : _GEN_11010; // @[icache.scala 138:25]
  wire [184:0] _GEN_15107 = lookup & dirty ? _GEN_14083 : _GEN_11011; // @[icache.scala 138:25]
  wire [184:0] _GEN_15108 = lookup & dirty ? _GEN_14084 : _GEN_11012; // @[icache.scala 138:25]
  wire [184:0] _GEN_15109 = lookup & dirty ? _GEN_14085 : _GEN_11013; // @[icache.scala 138:25]
  wire [184:0] _GEN_15110 = lookup & dirty ? _GEN_14086 : _GEN_11014; // @[icache.scala 138:25]
  wire [184:0] _GEN_15111 = lookup & dirty ? _GEN_14087 : _GEN_11015; // @[icache.scala 138:25]
  wire [184:0] _GEN_15112 = lookup & dirty ? _GEN_14088 : _GEN_11016; // @[icache.scala 138:25]
  wire [184:0] _GEN_15113 = lookup & dirty ? _GEN_14089 : _GEN_11017; // @[icache.scala 138:25]
  wire [184:0] _GEN_15114 = lookup & dirty ? _GEN_14090 : _GEN_11018; // @[icache.scala 138:25]
  wire [184:0] _GEN_15115 = lookup & dirty ? _GEN_14091 : _GEN_11019; // @[icache.scala 138:25]
  wire [184:0] _GEN_15116 = lookup & dirty ? _GEN_14092 : _GEN_11020; // @[icache.scala 138:25]
  wire [184:0] _GEN_15117 = lookup & dirty ? _GEN_14093 : _GEN_11021; // @[icache.scala 138:25]
  wire [184:0] _GEN_15118 = lookup & dirty ? _GEN_14094 : _GEN_11022; // @[icache.scala 138:25]
  wire [184:0] _GEN_15119 = lookup & dirty ? _GEN_14095 : _GEN_11023; // @[icache.scala 138:25]
  wire [184:0] _GEN_15120 = lookup & dirty ? _GEN_14096 : _GEN_11024; // @[icache.scala 138:25]
  wire [184:0] _GEN_15121 = lookup & dirty ? _GEN_14097 : _GEN_11025; // @[icache.scala 138:25]
  wire [184:0] _GEN_15122 = lookup & dirty ? _GEN_14098 : _GEN_11026; // @[icache.scala 138:25]
  wire [184:0] _GEN_15123 = lookup & dirty ? _GEN_14099 : _GEN_11027; // @[icache.scala 138:25]
  wire [184:0] _GEN_15124 = lookup & dirty ? _GEN_14100 : _GEN_11028; // @[icache.scala 138:25]
  wire [184:0] _GEN_15125 = lookup & dirty ? _GEN_14101 : _GEN_11029; // @[icache.scala 138:25]
  wire [184:0] _GEN_15126 = lookup & dirty ? _GEN_14102 : _GEN_11030; // @[icache.scala 138:25]
  wire [184:0] _GEN_15127 = lookup & dirty ? _GEN_14103 : _GEN_11031; // @[icache.scala 138:25]
  wire [184:0] _GEN_15128 = lookup & dirty ? _GEN_14104 : _GEN_11032; // @[icache.scala 138:25]
  wire [184:0] _GEN_15129 = lookup & dirty ? _GEN_14105 : _GEN_11033; // @[icache.scala 138:25]
  wire [184:0] _GEN_15130 = lookup & dirty ? _GEN_14106 : _GEN_11034; // @[icache.scala 138:25]
  wire [184:0] _GEN_15131 = lookup & dirty ? _GEN_14107 : _GEN_11035; // @[icache.scala 138:25]
  wire [184:0] _GEN_15132 = lookup & dirty ? _GEN_14108 : _GEN_11036; // @[icache.scala 138:25]
  wire [184:0] _GEN_15133 = lookup & dirty ? _GEN_14109 : _GEN_11037; // @[icache.scala 138:25]
  wire [184:0] _GEN_15134 = lookup & dirty ? _GEN_14110 : _GEN_11038; // @[icache.scala 138:25]
  wire [184:0] _GEN_15135 = lookup & dirty ? _GEN_14111 : _GEN_11039; // @[icache.scala 138:25]
  wire [184:0] _GEN_15136 = lookup & dirty ? _GEN_14112 : _GEN_11040; // @[icache.scala 138:25]
  wire [184:0] _GEN_15137 = lookup & dirty ? _GEN_14113 : _GEN_11041; // @[icache.scala 138:25]
  wire [184:0] _GEN_15138 = lookup & dirty ? _GEN_14114 : _GEN_11042; // @[icache.scala 138:25]
  wire [184:0] _GEN_15139 = lookup & dirty ? _GEN_14115 : _GEN_11043; // @[icache.scala 138:25]
  wire [184:0] _GEN_15140 = lookup & dirty ? _GEN_14116 : _GEN_11044; // @[icache.scala 138:25]
  wire [184:0] _GEN_15141 = lookup & dirty ? _GEN_14117 : _GEN_11045; // @[icache.scala 138:25]
  wire [184:0] _GEN_15142 = lookup & dirty ? _GEN_14118 : _GEN_11046; // @[icache.scala 138:25]
  wire [184:0] _GEN_15143 = lookup & dirty ? _GEN_14119 : _GEN_11047; // @[icache.scala 138:25]
  wire [184:0] _GEN_15144 = lookup & dirty ? _GEN_14120 : _GEN_11048; // @[icache.scala 138:25]
  wire [184:0] _GEN_15145 = lookup & dirty ? _GEN_14121 : _GEN_11049; // @[icache.scala 138:25]
  wire [184:0] _GEN_15146 = lookup & dirty ? _GEN_14122 : _GEN_11050; // @[icache.scala 138:25]
  wire [184:0] _GEN_15147 = lookup & dirty ? _GEN_14123 : _GEN_11051; // @[icache.scala 138:25]
  wire [184:0] _GEN_15148 = lookup & dirty ? _GEN_14124 : _GEN_11052; // @[icache.scala 138:25]
  wire [184:0] _GEN_15149 = lookup & dirty ? _GEN_14125 : _GEN_11053; // @[icache.scala 138:25]
  wire [184:0] _GEN_15150 = lookup & dirty ? _GEN_14126 : _GEN_11054; // @[icache.scala 138:25]
  wire [184:0] _GEN_15151 = lookup & dirty ? _GEN_14127 : _GEN_11055; // @[icache.scala 138:25]
  wire [184:0] _GEN_15152 = lookup & dirty ? _GEN_14128 : _GEN_11056; // @[icache.scala 138:25]
  wire [184:0] _GEN_15153 = lookup & dirty ? _GEN_14129 : _GEN_11057; // @[icache.scala 138:25]
  wire [184:0] _GEN_15154 = lookup & dirty ? _GEN_14130 : _GEN_11058; // @[icache.scala 138:25]
  wire [184:0] _GEN_15155 = lookup & dirty ? _GEN_14131 : _GEN_11059; // @[icache.scala 138:25]
  wire [184:0] _GEN_15156 = lookup & dirty ? _GEN_14132 : _GEN_11060; // @[icache.scala 138:25]
  wire [184:0] _GEN_15157 = lookup & dirty ? _GEN_14133 : _GEN_11061; // @[icache.scala 138:25]
  wire [184:0] _GEN_15158 = lookup & dirty ? _GEN_14134 : _GEN_11062; // @[icache.scala 138:25]
  wire [184:0] _GEN_15159 = lookup & dirty ? _GEN_14135 : _GEN_11063; // @[icache.scala 138:25]
  wire [184:0] _GEN_15160 = lookup & dirty ? _GEN_14136 : _GEN_11064; // @[icache.scala 138:25]
  wire [184:0] _GEN_15161 = lookup & dirty ? _GEN_14137 : _GEN_11065; // @[icache.scala 138:25]
  wire [184:0] _GEN_15162 = lookup & dirty ? _GEN_14138 : _GEN_11066; // @[icache.scala 138:25]
  wire [184:0] _GEN_15163 = lookup & dirty ? _GEN_14139 : _GEN_11067; // @[icache.scala 138:25]
  wire [184:0] _GEN_15164 = lookup & dirty ? _GEN_14140 : _GEN_11068; // @[icache.scala 138:25]
  wire [184:0] _GEN_15165 = lookup & dirty ? _GEN_14141 : _GEN_11069; // @[icache.scala 138:25]
  wire [184:0] _GEN_15166 = lookup & dirty ? _GEN_14142 : _GEN_11070; // @[icache.scala 138:25]
  wire [184:0] _GEN_15167 = lookup & dirty ? _GEN_14143 : _GEN_11071; // @[icache.scala 138:25]
  wire [184:0] _GEN_15168 = lookup & dirty ? _GEN_14144 : _GEN_11072; // @[icache.scala 138:25]
  wire [184:0] _GEN_15169 = lookup & dirty ? _GEN_14145 : _GEN_11073; // @[icache.scala 138:25]
  wire [184:0] _GEN_15170 = lookup & dirty ? _GEN_14146 : _GEN_11074; // @[icache.scala 138:25]
  wire [184:0] _GEN_15171 = lookup & dirty ? _GEN_14147 : _GEN_11075; // @[icache.scala 138:25]
  wire [184:0] _GEN_15172 = lookup & dirty ? _GEN_14148 : _GEN_11076; // @[icache.scala 138:25]
  wire [184:0] _GEN_15173 = lookup & dirty ? _GEN_14149 : _GEN_11077; // @[icache.scala 138:25]
  wire [184:0] _GEN_15174 = lookup & dirty ? _GEN_14150 : _GEN_11078; // @[icache.scala 138:25]
  wire [184:0] _GEN_15175 = lookup & dirty ? _GEN_14151 : _GEN_11079; // @[icache.scala 138:25]
  wire [184:0] _GEN_15176 = lookup & dirty ? _GEN_14152 : _GEN_11080; // @[icache.scala 138:25]
  wire [184:0] _GEN_15177 = lookup & dirty ? _GEN_14153 : _GEN_11081; // @[icache.scala 138:25]
  wire [184:0] _GEN_15178 = lookup & dirty ? _GEN_14154 : _GEN_11082; // @[icache.scala 138:25]
  wire [184:0] _GEN_15179 = lookup & dirty ? _GEN_14155 : _GEN_11083; // @[icache.scala 138:25]
  wire [184:0] _GEN_15180 = lookup & dirty ? _GEN_14156 : _GEN_11084; // @[icache.scala 138:25]
  wire [184:0] _GEN_15181 = lookup & dirty ? _GEN_14157 : _GEN_11085; // @[icache.scala 138:25]
  wire [184:0] _GEN_15182 = lookup & dirty ? _GEN_14158 : _GEN_11086; // @[icache.scala 138:25]
  wire [184:0] _GEN_15183 = lookup & dirty ? _GEN_14159 : _GEN_11087; // @[icache.scala 138:25]
  wire [184:0] _GEN_15184 = lookup & dirty ? _GEN_14160 : _GEN_11088; // @[icache.scala 138:25]
  wire [184:0] _GEN_15185 = lookup & dirty ? _GEN_14161 : _GEN_11089; // @[icache.scala 138:25]
  wire [184:0] _GEN_15186 = lookup & dirty ? _GEN_14162 : _GEN_11090; // @[icache.scala 138:25]
  wire [184:0] _GEN_15187 = lookup & dirty ? _GEN_14163 : _GEN_11091; // @[icache.scala 138:25]
  wire [184:0] _GEN_15188 = lookup & dirty ? _GEN_14164 : _GEN_11092; // @[icache.scala 138:25]
  wire [184:0] _GEN_15189 = lookup & dirty ? _GEN_14165 : _GEN_11093; // @[icache.scala 138:25]
  wire [184:0] _GEN_15190 = lookup & dirty ? _GEN_14166 : _GEN_11094; // @[icache.scala 138:25]
  wire [184:0] _GEN_15191 = lookup & dirty ? _GEN_14167 : _GEN_11095; // @[icache.scala 138:25]
  wire [184:0] _GEN_15192 = lookup & dirty ? _GEN_14168 : _GEN_11096; // @[icache.scala 138:25]
  wire [184:0] _GEN_15193 = lookup & dirty ? _GEN_14169 : _GEN_11097; // @[icache.scala 138:25]
  wire [184:0] _GEN_15194 = lookup & dirty ? _GEN_14170 : _GEN_11098; // @[icache.scala 138:25]
  wire [184:0] _GEN_15195 = lookup & dirty ? _GEN_14171 : _GEN_11099; // @[icache.scala 138:25]
  wire [184:0] _GEN_15196 = lookup & dirty ? _GEN_14172 : _GEN_11100; // @[icache.scala 138:25]
  wire [184:0] _GEN_15197 = lookup & dirty ? _GEN_14173 : _GEN_11101; // @[icache.scala 138:25]
  wire [184:0] _GEN_15198 = lookup & dirty ? _GEN_14174 : _GEN_11102; // @[icache.scala 138:25]
  wire [184:0] _GEN_15199 = lookup & dirty ? _GEN_14175 : _GEN_11103; // @[icache.scala 138:25]
  wire [184:0] _GEN_15200 = lookup & dirty ? _GEN_14176 : _GEN_11104; // @[icache.scala 138:25]
  wire [184:0] _GEN_15201 = lookup & dirty ? _GEN_14177 : _GEN_11105; // @[icache.scala 138:25]
  wire [184:0] _GEN_15202 = lookup & dirty ? _GEN_14178 : _GEN_11106; // @[icache.scala 138:25]
  wire [184:0] _GEN_15203 = lookup & dirty ? _GEN_14179 : _GEN_11107; // @[icache.scala 138:25]
  wire [184:0] _GEN_15204 = lookup & dirty ? _GEN_14180 : _GEN_11108; // @[icache.scala 138:25]
  wire [184:0] _GEN_15205 = lookup & dirty ? _GEN_14181 : _GEN_11109; // @[icache.scala 138:25]
  wire [184:0] _GEN_15206 = lookup & dirty ? _GEN_14182 : _GEN_11110; // @[icache.scala 138:25]
  wire [184:0] _GEN_15207 = lookup & dirty ? _GEN_14183 : _GEN_11111; // @[icache.scala 138:25]
  wire [184:0] _GEN_15208 = lookup & dirty ? _GEN_14184 : _GEN_11112; // @[icache.scala 138:25]
  wire [184:0] _GEN_15209 = lookup & dirty ? _GEN_14185 : _GEN_11113; // @[icache.scala 138:25]
  wire [184:0] _GEN_15210 = lookup & dirty ? _GEN_14186 : _GEN_11114; // @[icache.scala 138:25]
  wire [184:0] _GEN_15211 = lookup & dirty ? _GEN_14187 : _GEN_11115; // @[icache.scala 138:25]
  wire [184:0] _GEN_15212 = lookup & dirty ? _GEN_14188 : _GEN_11116; // @[icache.scala 138:25]
  wire [184:0] _GEN_15213 = lookup & dirty ? _GEN_14189 : _GEN_11117; // @[icache.scala 138:25]
  wire [184:0] _GEN_15214 = lookup & dirty ? _GEN_14190 : _GEN_11118; // @[icache.scala 138:25]
  wire [184:0] _GEN_15215 = lookup & dirty ? _GEN_14191 : _GEN_11119; // @[icache.scala 138:25]
  wire [184:0] _GEN_15216 = lookup & dirty ? _GEN_14192 : _GEN_11120; // @[icache.scala 138:25]
  wire [184:0] _GEN_15217 = lookup & dirty ? _GEN_14193 : _GEN_11121; // @[icache.scala 138:25]
  wire [184:0] _GEN_15218 = lookup & dirty ? _GEN_14194 : _GEN_11122; // @[icache.scala 138:25]
  wire [184:0] _GEN_15219 = lookup & dirty ? _GEN_14195 : _GEN_11123; // @[icache.scala 138:25]
  wire [184:0] _GEN_15220 = lookup & dirty ? _GEN_14196 : _GEN_11124; // @[icache.scala 138:25]
  wire [184:0] _GEN_15221 = lookup & dirty ? _GEN_14197 : _GEN_11125; // @[icache.scala 138:25]
  wire [184:0] _GEN_15222 = lookup & dirty ? _GEN_14198 : _GEN_11126; // @[icache.scala 138:25]
  wire [184:0] _GEN_15223 = lookup & dirty ? _GEN_14199 : _GEN_11127; // @[icache.scala 138:25]
  wire [184:0] _GEN_15224 = lookup & dirty ? _GEN_14200 : _GEN_11128; // @[icache.scala 138:25]
  wire [184:0] _GEN_15225 = lookup & dirty ? _GEN_14201 : _GEN_11129; // @[icache.scala 138:25]
  wire [184:0] _GEN_15226 = lookup & dirty ? _GEN_14202 : _GEN_11130; // @[icache.scala 138:25]
  wire [184:0] _GEN_15227 = lookup & dirty ? _GEN_14203 : _GEN_11131; // @[icache.scala 138:25]
  wire [184:0] _GEN_15228 = lookup & dirty ? _GEN_14204 : _GEN_11132; // @[icache.scala 138:25]
  wire [184:0] _GEN_15229 = lookup & dirty ? _GEN_14205 : _GEN_11133; // @[icache.scala 138:25]
  wire [184:0] _GEN_15230 = lookup & dirty ? _GEN_14206 : _GEN_11134; // @[icache.scala 138:25]
  wire [184:0] _GEN_15231 = lookup & dirty ? _GEN_14207 : _GEN_11135; // @[icache.scala 138:25]
  wire [184:0] _GEN_15232 = lookup & dirty ? _GEN_14208 : _GEN_11136; // @[icache.scala 138:25]
  wire [184:0] _GEN_15233 = lookup & dirty ? _GEN_14209 : _GEN_11137; // @[icache.scala 138:25]
  wire [184:0] _GEN_15234 = lookup & dirty ? _GEN_14210 : _GEN_11138; // @[icache.scala 138:25]
  wire [184:0] _GEN_15235 = lookup & dirty ? _GEN_14211 : _GEN_11139; // @[icache.scala 138:25]
  wire [184:0] _GEN_15236 = lookup & dirty ? _GEN_14212 : _GEN_11140; // @[icache.scala 138:25]
  wire [184:0] _GEN_15237 = lookup & dirty ? _GEN_14213 : _GEN_11141; // @[icache.scala 138:25]
  wire [184:0] _GEN_15238 = lookup & dirty ? _GEN_14214 : _GEN_11142; // @[icache.scala 138:25]
  wire [184:0] _GEN_15239 = lookup & dirty ? _GEN_14215 : _GEN_11143; // @[icache.scala 138:25]
  wire [184:0] _GEN_15240 = lookup & dirty ? _GEN_14216 : _GEN_11144; // @[icache.scala 138:25]
  wire [184:0] _GEN_15241 = lookup & dirty ? _GEN_14217 : _GEN_11145; // @[icache.scala 138:25]
  wire [184:0] _GEN_15242 = lookup & dirty ? _GEN_14218 : _GEN_11146; // @[icache.scala 138:25]
  wire [184:0] _GEN_15243 = lookup & dirty ? _GEN_14219 : _GEN_11147; // @[icache.scala 138:25]
  wire [184:0] _GEN_15244 = lookup & dirty ? _GEN_14220 : _GEN_11148; // @[icache.scala 138:25]
  wire [184:0] _GEN_15245 = lookup & dirty ? _GEN_14221 : _GEN_11149; // @[icache.scala 138:25]
  wire [184:0] _GEN_15246 = lookup & dirty ? _GEN_14222 : _GEN_11150; // @[icache.scala 138:25]
  wire [184:0] _GEN_15247 = lookup & dirty ? _GEN_14223 : _GEN_11151; // @[icache.scala 138:25]
  wire [184:0] _GEN_15248 = lookup & dirty ? _GEN_14224 : _GEN_11152; // @[icache.scala 138:25]
  wire [184:0] _GEN_15249 = lookup & dirty ? _GEN_14225 : _GEN_11153; // @[icache.scala 138:25]
  wire [184:0] _GEN_15250 = lookup & dirty ? _GEN_14226 : _GEN_11154; // @[icache.scala 138:25]
  wire [184:0] _GEN_15251 = lookup & dirty ? _GEN_14227 : _GEN_11155; // @[icache.scala 138:25]
  wire [184:0] _GEN_15252 = lookup & dirty ? _GEN_14228 : _GEN_11156; // @[icache.scala 138:25]
  wire [184:0] _GEN_15253 = lookup & dirty ? _GEN_14229 : _GEN_11157; // @[icache.scala 138:25]
  wire [184:0] _GEN_15254 = lookup & dirty ? _GEN_14230 : _GEN_11158; // @[icache.scala 138:25]
  wire [184:0] _GEN_15255 = lookup & dirty ? _GEN_14231 : _GEN_11159; // @[icache.scala 138:25]
  wire [184:0] _GEN_15256 = lookup & dirty ? _GEN_14232 : _GEN_11160; // @[icache.scala 138:25]
  wire [184:0] _GEN_15257 = lookup & dirty ? _GEN_14233 : _GEN_11161; // @[icache.scala 138:25]
  wire [184:0] _GEN_15258 = lookup & dirty ? _GEN_14234 : _GEN_11162; // @[icache.scala 138:25]
  wire [184:0] _GEN_15259 = lookup & dirty ? _GEN_14235 : _GEN_11163; // @[icache.scala 138:25]
  wire [184:0] _GEN_15260 = lookup & dirty ? _GEN_14236 : _GEN_11164; // @[icache.scala 138:25]
  wire [184:0] _GEN_15261 = lookup & dirty ? _GEN_14237 : _GEN_11165; // @[icache.scala 138:25]
  wire [184:0] _GEN_15262 = lookup & dirty ? _GEN_14238 : _GEN_11166; // @[icache.scala 138:25]
  wire [184:0] _GEN_15263 = lookup & dirty ? _GEN_14239 : _GEN_11167; // @[icache.scala 138:25]
  wire [184:0] _GEN_15264 = lookup & dirty ? _GEN_14240 : _GEN_11168; // @[icache.scala 138:25]
  wire [184:0] _GEN_15265 = lookup & dirty ? _GEN_14241 : _GEN_11169; // @[icache.scala 138:25]
  wire [184:0] _GEN_15266 = lookup & dirty ? _GEN_14242 : _GEN_11170; // @[icache.scala 138:25]
  wire [184:0] _GEN_15267 = lookup & dirty ? _GEN_14243 : _GEN_11171; // @[icache.scala 138:25]
  wire [184:0] _GEN_15268 = lookup & dirty ? _GEN_14244 : _GEN_11172; // @[icache.scala 138:25]
  wire [184:0] _GEN_15269 = lookup & dirty ? _GEN_14245 : _GEN_11173; // @[icache.scala 138:25]
  wire [184:0] _GEN_15270 = lookup & dirty ? _GEN_14246 : _GEN_11174; // @[icache.scala 138:25]
  wire [184:0] _GEN_15271 = lookup & dirty ? _GEN_14247 : _GEN_11175; // @[icache.scala 138:25]
  wire [184:0] _GEN_15272 = lookup & dirty ? _GEN_14248 : _GEN_11176; // @[icache.scala 138:25]
  wire [184:0] _GEN_15273 = lookup & dirty ? _GEN_14249 : _GEN_11177; // @[icache.scala 138:25]
  wire [184:0] _GEN_15274 = lookup & dirty ? _GEN_14250 : _GEN_11178; // @[icache.scala 138:25]
  wire [184:0] _GEN_15275 = lookup & dirty ? _GEN_14251 : _GEN_11179; // @[icache.scala 138:25]
  wire [184:0] _GEN_15276 = lookup & dirty ? _GEN_14252 : _GEN_11180; // @[icache.scala 138:25]
  wire [184:0] _GEN_15277 = lookup & dirty ? _GEN_14253 : _GEN_11181; // @[icache.scala 138:25]
  wire [184:0] _GEN_15278 = lookup & dirty ? _GEN_14254 : _GEN_11182; // @[icache.scala 138:25]
  wire [184:0] _GEN_15279 = lookup & dirty ? _GEN_14255 : _GEN_11183; // @[icache.scala 138:25]
  wire [184:0] _GEN_15280 = lookup & dirty ? _GEN_14256 : _GEN_11184; // @[icache.scala 138:25]
  wire [184:0] _GEN_15281 = lookup & dirty ? _GEN_14257 : _GEN_11185; // @[icache.scala 138:25]
  wire [184:0] _GEN_15282 = lookup & dirty ? _GEN_14258 : _GEN_11186; // @[icache.scala 138:25]
  wire [184:0] _GEN_15283 = lookup & dirty ? _GEN_14259 : _GEN_11187; // @[icache.scala 138:25]
  wire [184:0] _GEN_15284 = lookup & dirty ? _GEN_14260 : _GEN_11188; // @[icache.scala 138:25]
  wire [184:0] _GEN_15285 = lookup & dirty ? _GEN_14261 : _GEN_11189; // @[icache.scala 138:25]
  wire [184:0] _GEN_15286 = lookup & dirty ? _GEN_14262 : _GEN_11190; // @[icache.scala 138:25]
  wire [184:0] _GEN_15287 = lookup & dirty ? _GEN_14263 : _GEN_11191; // @[icache.scala 138:25]
  wire [184:0] _GEN_15288 = lookup & dirty ? _GEN_14264 : _GEN_11192; // @[icache.scala 138:25]
  wire [184:0] _GEN_15289 = lookup & dirty ? _GEN_14265 : _GEN_11193; // @[icache.scala 138:25]
  wire [184:0] _GEN_15290 = lookup & dirty ? _GEN_14266 : _GEN_11194; // @[icache.scala 138:25]
  wire [184:0] _GEN_15291 = lookup & dirty ? _GEN_14267 : _GEN_11195; // @[icache.scala 138:25]
  wire [184:0] _GEN_15292 = lookup & dirty ? _GEN_14268 : _GEN_11196; // @[icache.scala 138:25]
  wire [184:0] _GEN_15293 = lookup & dirty ? _GEN_14269 : _GEN_11197; // @[icache.scala 138:25]
  wire [184:0] _GEN_15294 = lookup & dirty ? _GEN_14270 : _GEN_11198; // @[icache.scala 138:25]
  wire [184:0] _GEN_15295 = lookup & dirty ? _GEN_14271 : _GEN_11199; // @[icache.scala 138:25]
  wire [184:0] _GEN_15296 = lookup & dirty ? _GEN_14272 : _GEN_11200; // @[icache.scala 138:25]
  wire [184:0] _GEN_15297 = lookup & dirty ? _GEN_14273 : _GEN_11201; // @[icache.scala 138:25]
  wire [184:0] _GEN_15298 = lookup & dirty ? _GEN_14274 : _GEN_11202; // @[icache.scala 138:25]
  wire [184:0] _GEN_15299 = lookup & dirty ? _GEN_14275 : _GEN_11203; // @[icache.scala 138:25]
  wire [184:0] _GEN_15300 = lookup & dirty ? _GEN_14276 : _GEN_11204; // @[icache.scala 138:25]
  wire [184:0] _GEN_15301 = lookup & dirty ? _GEN_14277 : _GEN_11205; // @[icache.scala 138:25]
  wire [184:0] _GEN_15302 = lookup & dirty ? _GEN_14278 : _GEN_11206; // @[icache.scala 138:25]
  wire [184:0] _GEN_15303 = lookup & dirty ? _GEN_14279 : _GEN_11207; // @[icache.scala 138:25]
  wire [184:0] _GEN_15304 = lookup & dirty ? _GEN_14280 : _GEN_11208; // @[icache.scala 138:25]
  wire [184:0] _GEN_15305 = lookup & dirty ? _GEN_14281 : _GEN_11209; // @[icache.scala 138:25]
  wire [184:0] _GEN_15306 = lookup & dirty ? _GEN_14282 : _GEN_11210; // @[icache.scala 138:25]
  wire [184:0] _GEN_15307 = lookup & dirty ? _GEN_14283 : _GEN_11211; // @[icache.scala 138:25]
  wire [184:0] _GEN_15308 = lookup & dirty ? _GEN_14284 : _GEN_11212; // @[icache.scala 138:25]
  wire [184:0] _GEN_15309 = lookup & dirty ? _GEN_14285 : _GEN_11213; // @[icache.scala 138:25]
  wire [184:0] _GEN_15310 = lookup & dirty ? _GEN_14286 : _GEN_11214; // @[icache.scala 138:25]
  wire [184:0] _GEN_15311 = lookup & dirty ? _GEN_14287 : _GEN_11215; // @[icache.scala 138:25]
  wire [184:0] _GEN_15312 = lookup & dirty ? _GEN_14288 : _GEN_11216; // @[icache.scala 138:25]
  wire [184:0] _GEN_15313 = lookup & dirty ? _GEN_14289 : _GEN_11217; // @[icache.scala 138:25]
  wire [184:0] _GEN_15314 = lookup & dirty ? _GEN_14290 : _GEN_11218; // @[icache.scala 138:25]
  wire [184:0] _GEN_15315 = lookup & dirty ? _GEN_14291 : _GEN_11219; // @[icache.scala 138:25]
  wire [184:0] _GEN_15316 = lookup & dirty ? _GEN_14292 : _GEN_11220; // @[icache.scala 138:25]
  wire [184:0] _GEN_15317 = lookup & dirty ? _GEN_14293 : _GEN_11221; // @[icache.scala 138:25]
  wire [184:0] _GEN_15318 = lookup & dirty ? _GEN_14294 : _GEN_11222; // @[icache.scala 138:25]
  wire [184:0] _GEN_15319 = lookup & dirty ? _GEN_14295 : _GEN_11223; // @[icache.scala 138:25]
  wire [184:0] _GEN_15320 = lookup & dirty ? _GEN_14296 : _GEN_11224; // @[icache.scala 138:25]
  wire [184:0] _GEN_15321 = lookup & dirty ? _GEN_14297 : _GEN_11225; // @[icache.scala 138:25]
  wire [184:0] _GEN_15322 = lookup & dirty ? _GEN_14298 : _GEN_11226; // @[icache.scala 138:25]
  wire [184:0] _GEN_15323 = lookup & dirty ? _GEN_14299 : _GEN_11227; // @[icache.scala 138:25]
  wire [184:0] _GEN_15324 = lookup & dirty ? _GEN_14300 : _GEN_11228; // @[icache.scala 138:25]
  wire [184:0] _GEN_15325 = lookup & dirty ? _GEN_14301 : _GEN_11229; // @[icache.scala 138:25]
  wire [184:0] _GEN_15326 = lookup & dirty ? _GEN_14302 : _GEN_11230; // @[icache.scala 138:25]
  wire [184:0] _GEN_15327 = lookup & dirty ? _GEN_14303 : _GEN_11231; // @[icache.scala 138:25]
  wire [184:0] _GEN_15328 = lookup & dirty ? _GEN_14304 : _GEN_11232; // @[icache.scala 138:25]
  wire [184:0] _GEN_15329 = lookup & dirty ? _GEN_14305 : _GEN_11233; // @[icache.scala 138:25]
  wire [184:0] _GEN_15330 = lookup & dirty ? _GEN_14306 : _GEN_11234; // @[icache.scala 138:25]
  wire [184:0] _GEN_15331 = lookup & dirty ? _GEN_14307 : _GEN_11235; // @[icache.scala 138:25]
  wire [184:0] _GEN_15332 = lookup & dirty ? _GEN_14308 : _GEN_11236; // @[icache.scala 138:25]
  wire [184:0] _GEN_15333 = lookup & dirty ? _GEN_14309 : _GEN_11237; // @[icache.scala 138:25]
  wire [184:0] _GEN_15334 = lookup & dirty ? _GEN_14310 : _GEN_11238; // @[icache.scala 138:25]
  wire [184:0] _GEN_15335 = lookup & dirty ? _GEN_14311 : _GEN_11239; // @[icache.scala 138:25]
  wire [184:0] _GEN_15336 = lookup & dirty ? _GEN_14312 : _GEN_11240; // @[icache.scala 138:25]
  wire [184:0] _GEN_15337 = lookup & dirty ? _GEN_14313 : _GEN_11241; // @[icache.scala 138:25]
  wire [184:0] _GEN_15338 = lookup & dirty ? _GEN_14314 : _GEN_11242; // @[icache.scala 138:25]
  wire [184:0] _GEN_15339 = lookup & dirty ? _GEN_14315 : _GEN_11243; // @[icache.scala 138:25]
  wire [184:0] _GEN_15340 = lookup & dirty ? _GEN_14316 : _GEN_11244; // @[icache.scala 138:25]
  wire [184:0] _GEN_15341 = lookup & dirty ? _GEN_14317 : _GEN_11245; // @[icache.scala 138:25]
  wire [184:0] _GEN_15342 = lookup & dirty ? _GEN_14318 : _GEN_11246; // @[icache.scala 138:25]
  wire [184:0] _GEN_15343 = lookup & dirty ? _GEN_14319 : _GEN_11247; // @[icache.scala 138:25]
  wire [184:0] _GEN_15344 = lookup & dirty ? _GEN_14320 : _GEN_11248; // @[icache.scala 138:25]
  wire [184:0] _GEN_15345 = lookup & dirty ? _GEN_14321 : _GEN_11249; // @[icache.scala 138:25]
  wire [184:0] _GEN_15346 = lookup & dirty ? _GEN_14322 : _GEN_11250; // @[icache.scala 138:25]
  wire [184:0] _GEN_15347 = lookup & dirty ? _GEN_14323 : _GEN_11251; // @[icache.scala 138:25]
  wire [184:0] _GEN_15348 = lookup & dirty ? _GEN_14324 : _GEN_11252; // @[icache.scala 138:25]
  wire [184:0] _GEN_15349 = lookup & dirty ? _GEN_14325 : _GEN_11253; // @[icache.scala 138:25]
  wire [184:0] _GEN_15350 = lookup & dirty ? _GEN_14326 : _GEN_11254; // @[icache.scala 138:25]
  wire [184:0] _GEN_15351 = lookup & dirty ? _GEN_14327 : _GEN_11255; // @[icache.scala 138:25]
  wire [184:0] _GEN_15352 = lookup & dirty ? _GEN_14328 : _GEN_11256; // @[icache.scala 138:25]
  wire [184:0] _GEN_15353 = lookup & dirty ? _GEN_14329 : _GEN_11257; // @[icache.scala 138:25]
  wire [184:0] _GEN_15354 = lookup & dirty ? _GEN_14330 : _GEN_11258; // @[icache.scala 138:25]
  wire [184:0] _GEN_15355 = lookup & dirty ? _GEN_14331 : _GEN_11259; // @[icache.scala 138:25]
  wire [184:0] _GEN_15356 = lookup & dirty ? _GEN_14332 : _GEN_11260; // @[icache.scala 138:25]
  wire [184:0] _GEN_15357 = lookup & dirty ? _GEN_14333 : _GEN_11261; // @[icache.scala 138:25]
  wire [184:0] _GEN_15358 = lookup & dirty ? _GEN_14334 : _GEN_11262; // @[icache.scala 138:25]
  wire [184:0] _GEN_15359 = lookup & dirty ? _GEN_14335 : _GEN_11263; // @[icache.scala 138:25]
  wire [184:0] _GEN_15360 = lookup & dirty ? _GEN_14336 : _GEN_11264; // @[icache.scala 138:25]
  wire [184:0] _GEN_15361 = lookup & dirty ? _GEN_14337 : _GEN_11265; // @[icache.scala 138:25]
  wire [184:0] _GEN_15362 = lookup & dirty ? _GEN_14338 : _GEN_11266; // @[icache.scala 138:25]
  wire [184:0] _GEN_15363 = lookup & dirty ? _GEN_14339 : _GEN_11267; // @[icache.scala 138:25]
  wire [184:0] _GEN_15364 = lookup & dirty ? _GEN_14340 : _GEN_11268; // @[icache.scala 138:25]
  wire [184:0] _GEN_15365 = lookup & dirty ? _GEN_14341 : _GEN_11269; // @[icache.scala 138:25]
  wire [184:0] _GEN_15366 = lookup & dirty ? _GEN_14342 : _GEN_11270; // @[icache.scala 138:25]
  wire [184:0] _GEN_15367 = lookup & dirty ? _GEN_14343 : _GEN_11271; // @[icache.scala 138:25]
  wire [184:0] _GEN_15368 = lookup & dirty ? _GEN_14344 : _GEN_11272; // @[icache.scala 138:25]
  wire [184:0] _GEN_15369 = lookup & dirty ? _GEN_14345 : _GEN_11273; // @[icache.scala 138:25]
  wire [184:0] _GEN_15370 = lookup & dirty ? _GEN_14346 : _GEN_11274; // @[icache.scala 138:25]
  wire [184:0] _GEN_15371 = lookup & dirty ? _GEN_14347 : _GEN_11275; // @[icache.scala 138:25]
  wire [184:0] _GEN_15372 = lookup & dirty ? _GEN_14348 : _GEN_11276; // @[icache.scala 138:25]
  wire [184:0] _GEN_15373 = lookup & dirty ? _GEN_14349 : _GEN_11277; // @[icache.scala 138:25]
  wire [184:0] _cache_data_T_17 = {1'h1,_GEN_4095[183],cpu_tag,io_rd_data}; // @[Cat.scala 31:58]
  assign io_rdata = reg_rdata; // @[icache.scala 164:19 165:14]
  assign io_addr_ok = lookup & hit; // @[icache.scala 157:24]
  assign io_data_ok = delay; // @[icache.scala 158:23]
  assign io_rd_req = state == 2'h3; // @[icache.scala 27:66]
  assign io_rd_addr = io_addr[31:0];
  always @(posedge clock) begin
    if (reset) begin // @[icache.scala 23:67]
      state <= 2'h0; // @[icache.scala 23:67]
    end else if (reset) begin // @[icache.scala 128:24]
      state <= 2'h0; // @[icache.scala 129:11]
    end else if (2'h0 == state) begin // @[icache.scala 53:17]
      if (io_valid) begin // @[icache.scala 55:22]
        state <= 2'h1; // @[icache.scala 56:15]
      end else begin
        state <= 2'h0; // @[icache.scala 58:15]
      end
    end else if (2'h1 == state) begin // @[icache.scala 53:17]
      state <= _GEN_4099;
    end else begin
      state <= _GEN_4103;
    end
    if (reset) begin // @[icache.scala 40:26]
      reg_rdata <= 64'h0; // @[icache.scala 40:26]
    end else if (_T_5 & way1_hit) begin // @[icache.scala 115:35]
      reg_rdata <= _GEN_2047[63:0]; // @[icache.scala 124:15]
    end else if (lookup & hit & way0_hit) begin // @[icache.scala 103:35]
      reg_rdata <= _GEN_1023[63:0]; // @[icache.scala 112:15]
    end
    if (reset) begin // @[icache.scala 41:25]
      delay <= 1'h0; // @[icache.scala 41:25]
    end else begin
      delay <= io_addr_ok;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_0 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_0 <= _GEN_14350;
      end
    end else begin
      cache_data_0 <= _GEN_14350;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1 <= _GEN_14351;
      end
    end else begin
      cache_data_1 <= _GEN_14351;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_2 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_2 <= _GEN_14352;
      end
    end else begin
      cache_data_2 <= _GEN_14352;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_3 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_3 <= _GEN_14353;
      end
    end else begin
      cache_data_3 <= _GEN_14353;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_4 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_4 <= _GEN_14354;
      end
    end else begin
      cache_data_4 <= _GEN_14354;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_5 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_5 <= _GEN_14355;
      end
    end else begin
      cache_data_5 <= _GEN_14355;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_6 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_6 <= _GEN_14356;
      end
    end else begin
      cache_data_6 <= _GEN_14356;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_7 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_7 <= _GEN_14357;
      end
    end else begin
      cache_data_7 <= _GEN_14357;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_8 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_8 <= _GEN_14358;
      end
    end else begin
      cache_data_8 <= _GEN_14358;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_9 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_9 <= _GEN_14359;
      end
    end else begin
      cache_data_9 <= _GEN_14359;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'ha == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_10 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_10 <= _GEN_14360;
      end
    end else begin
      cache_data_10 <= _GEN_14360;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_11 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_11 <= _GEN_14361;
      end
    end else begin
      cache_data_11 <= _GEN_14361;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_12 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_12 <= _GEN_14362;
      end
    end else begin
      cache_data_12 <= _GEN_14362;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_13 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_13 <= _GEN_14363;
      end
    end else begin
      cache_data_13 <= _GEN_14363;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'he == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_14 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_14 <= _GEN_14364;
      end
    end else begin
      cache_data_14 <= _GEN_14364;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hf == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_15 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_15 <= _GEN_14365;
      end
    end else begin
      cache_data_15 <= _GEN_14365;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h10 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_16 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_16 <= _GEN_14366;
      end
    end else begin
      cache_data_16 <= _GEN_14366;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h11 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_17 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_17 <= _GEN_14367;
      end
    end else begin
      cache_data_17 <= _GEN_14367;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h12 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_18 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_18 <= _GEN_14368;
      end
    end else begin
      cache_data_18 <= _GEN_14368;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h13 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_19 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_19 <= _GEN_14369;
      end
    end else begin
      cache_data_19 <= _GEN_14369;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h14 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_20 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_20 <= _GEN_14370;
      end
    end else begin
      cache_data_20 <= _GEN_14370;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h15 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_21 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_21 <= _GEN_14371;
      end
    end else begin
      cache_data_21 <= _GEN_14371;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h16 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_22 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_22 <= _GEN_14372;
      end
    end else begin
      cache_data_22 <= _GEN_14372;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h17 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_23 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_23 <= _GEN_14373;
      end
    end else begin
      cache_data_23 <= _GEN_14373;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h18 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_24 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_24 <= _GEN_14374;
      end
    end else begin
      cache_data_24 <= _GEN_14374;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h19 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_25 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_25 <= _GEN_14375;
      end
    end else begin
      cache_data_25 <= _GEN_14375;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_26 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_26 <= _GEN_14376;
      end
    end else begin
      cache_data_26 <= _GEN_14376;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_27 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_27 <= _GEN_14377;
      end
    end else begin
      cache_data_27 <= _GEN_14377;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_28 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_28 <= _GEN_14378;
      end
    end else begin
      cache_data_28 <= _GEN_14378;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_29 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_29 <= _GEN_14379;
      end
    end else begin
      cache_data_29 <= _GEN_14379;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_30 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_30 <= _GEN_14380;
      end
    end else begin
      cache_data_30 <= _GEN_14380;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_31 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_31 <= _GEN_14381;
      end
    end else begin
      cache_data_31 <= _GEN_14381;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h20 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_32 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_32 <= _GEN_14382;
      end
    end else begin
      cache_data_32 <= _GEN_14382;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h21 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_33 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_33 <= _GEN_14383;
      end
    end else begin
      cache_data_33 <= _GEN_14383;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h22 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_34 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_34 <= _GEN_14384;
      end
    end else begin
      cache_data_34 <= _GEN_14384;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h23 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_35 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_35 <= _GEN_14385;
      end
    end else begin
      cache_data_35 <= _GEN_14385;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h24 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_36 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_36 <= _GEN_14386;
      end
    end else begin
      cache_data_36 <= _GEN_14386;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h25 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_37 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_37 <= _GEN_14387;
      end
    end else begin
      cache_data_37 <= _GEN_14387;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h26 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_38 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_38 <= _GEN_14388;
      end
    end else begin
      cache_data_38 <= _GEN_14388;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h27 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_39 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_39 <= _GEN_14389;
      end
    end else begin
      cache_data_39 <= _GEN_14389;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h28 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_40 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_40 <= _GEN_14390;
      end
    end else begin
      cache_data_40 <= _GEN_14390;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h29 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_41 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_41 <= _GEN_14391;
      end
    end else begin
      cache_data_41 <= _GEN_14391;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_42 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_42 <= _GEN_14392;
      end
    end else begin
      cache_data_42 <= _GEN_14392;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_43 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_43 <= _GEN_14393;
      end
    end else begin
      cache_data_43 <= _GEN_14393;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_44 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_44 <= _GEN_14394;
      end
    end else begin
      cache_data_44 <= _GEN_14394;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_45 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_45 <= _GEN_14395;
      end
    end else begin
      cache_data_45 <= _GEN_14395;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_46 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_46 <= _GEN_14396;
      end
    end else begin
      cache_data_46 <= _GEN_14396;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_47 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_47 <= _GEN_14397;
      end
    end else begin
      cache_data_47 <= _GEN_14397;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h30 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_48 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_48 <= _GEN_14398;
      end
    end else begin
      cache_data_48 <= _GEN_14398;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h31 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_49 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_49 <= _GEN_14399;
      end
    end else begin
      cache_data_49 <= _GEN_14399;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h32 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_50 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_50 <= _GEN_14400;
      end
    end else begin
      cache_data_50 <= _GEN_14400;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h33 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_51 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_51 <= _GEN_14401;
      end
    end else begin
      cache_data_51 <= _GEN_14401;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h34 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_52 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_52 <= _GEN_14402;
      end
    end else begin
      cache_data_52 <= _GEN_14402;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h35 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_53 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_53 <= _GEN_14403;
      end
    end else begin
      cache_data_53 <= _GEN_14403;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h36 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_54 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_54 <= _GEN_14404;
      end
    end else begin
      cache_data_54 <= _GEN_14404;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h37 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_55 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_55 <= _GEN_14405;
      end
    end else begin
      cache_data_55 <= _GEN_14405;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h38 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_56 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_56 <= _GEN_14406;
      end
    end else begin
      cache_data_56 <= _GEN_14406;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h39 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_57 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_57 <= _GEN_14407;
      end
    end else begin
      cache_data_57 <= _GEN_14407;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_58 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_58 <= _GEN_14408;
      end
    end else begin
      cache_data_58 <= _GEN_14408;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_59 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_59 <= _GEN_14409;
      end
    end else begin
      cache_data_59 <= _GEN_14409;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_60 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_60 <= _GEN_14410;
      end
    end else begin
      cache_data_60 <= _GEN_14410;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_61 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_61 <= _GEN_14411;
      end
    end else begin
      cache_data_61 <= _GEN_14411;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_62 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_62 <= _GEN_14412;
      end
    end else begin
      cache_data_62 <= _GEN_14412;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_63 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_63 <= _GEN_14413;
      end
    end else begin
      cache_data_63 <= _GEN_14413;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h40 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_64 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_64 <= _GEN_14414;
      end
    end else begin
      cache_data_64 <= _GEN_14414;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h41 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_65 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_65 <= _GEN_14415;
      end
    end else begin
      cache_data_65 <= _GEN_14415;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h42 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_66 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_66 <= _GEN_14416;
      end
    end else begin
      cache_data_66 <= _GEN_14416;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h43 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_67 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_67 <= _GEN_14417;
      end
    end else begin
      cache_data_67 <= _GEN_14417;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h44 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_68 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_68 <= _GEN_14418;
      end
    end else begin
      cache_data_68 <= _GEN_14418;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h45 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_69 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_69 <= _GEN_14419;
      end
    end else begin
      cache_data_69 <= _GEN_14419;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h46 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_70 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_70 <= _GEN_14420;
      end
    end else begin
      cache_data_70 <= _GEN_14420;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h47 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_71 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_71 <= _GEN_14421;
      end
    end else begin
      cache_data_71 <= _GEN_14421;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h48 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_72 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_72 <= _GEN_14422;
      end
    end else begin
      cache_data_72 <= _GEN_14422;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h49 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_73 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_73 <= _GEN_14423;
      end
    end else begin
      cache_data_73 <= _GEN_14423;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h4a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_74 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_74 <= _GEN_14424;
      end
    end else begin
      cache_data_74 <= _GEN_14424;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h4b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_75 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_75 <= _GEN_14425;
      end
    end else begin
      cache_data_75 <= _GEN_14425;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h4c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_76 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_76 <= _GEN_14426;
      end
    end else begin
      cache_data_76 <= _GEN_14426;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h4d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_77 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_77 <= _GEN_14427;
      end
    end else begin
      cache_data_77 <= _GEN_14427;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h4e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_78 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_78 <= _GEN_14428;
      end
    end else begin
      cache_data_78 <= _GEN_14428;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h4f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_79 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_79 <= _GEN_14429;
      end
    end else begin
      cache_data_79 <= _GEN_14429;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h50 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_80 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_80 <= _GEN_14430;
      end
    end else begin
      cache_data_80 <= _GEN_14430;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h51 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_81 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_81 <= _GEN_14431;
      end
    end else begin
      cache_data_81 <= _GEN_14431;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h52 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_82 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_82 <= _GEN_14432;
      end
    end else begin
      cache_data_82 <= _GEN_14432;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h53 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_83 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_83 <= _GEN_14433;
      end
    end else begin
      cache_data_83 <= _GEN_14433;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h54 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_84 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_84 <= _GEN_14434;
      end
    end else begin
      cache_data_84 <= _GEN_14434;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h55 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_85 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_85 <= _GEN_14435;
      end
    end else begin
      cache_data_85 <= _GEN_14435;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h56 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_86 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_86 <= _GEN_14436;
      end
    end else begin
      cache_data_86 <= _GEN_14436;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h57 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_87 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_87 <= _GEN_14437;
      end
    end else begin
      cache_data_87 <= _GEN_14437;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h58 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_88 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_88 <= _GEN_14438;
      end
    end else begin
      cache_data_88 <= _GEN_14438;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h59 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_89 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_89 <= _GEN_14439;
      end
    end else begin
      cache_data_89 <= _GEN_14439;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h5a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_90 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_90 <= _GEN_14440;
      end
    end else begin
      cache_data_90 <= _GEN_14440;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h5b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_91 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_91 <= _GEN_14441;
      end
    end else begin
      cache_data_91 <= _GEN_14441;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h5c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_92 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_92 <= _GEN_14442;
      end
    end else begin
      cache_data_92 <= _GEN_14442;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h5d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_93 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_93 <= _GEN_14443;
      end
    end else begin
      cache_data_93 <= _GEN_14443;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h5e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_94 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_94 <= _GEN_14444;
      end
    end else begin
      cache_data_94 <= _GEN_14444;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h5f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_95 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_95 <= _GEN_14445;
      end
    end else begin
      cache_data_95 <= _GEN_14445;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h60 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_96 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_96 <= _GEN_14446;
      end
    end else begin
      cache_data_96 <= _GEN_14446;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h61 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_97 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_97 <= _GEN_14447;
      end
    end else begin
      cache_data_97 <= _GEN_14447;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h62 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_98 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_98 <= _GEN_14448;
      end
    end else begin
      cache_data_98 <= _GEN_14448;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h63 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_99 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_99 <= _GEN_14449;
      end
    end else begin
      cache_data_99 <= _GEN_14449;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h64 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_100 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_100 <= _GEN_14450;
      end
    end else begin
      cache_data_100 <= _GEN_14450;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h65 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_101 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_101 <= _GEN_14451;
      end
    end else begin
      cache_data_101 <= _GEN_14451;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h66 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_102 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_102 <= _GEN_14452;
      end
    end else begin
      cache_data_102 <= _GEN_14452;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h67 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_103 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_103 <= _GEN_14453;
      end
    end else begin
      cache_data_103 <= _GEN_14453;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h68 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_104 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_104 <= _GEN_14454;
      end
    end else begin
      cache_data_104 <= _GEN_14454;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h69 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_105 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_105 <= _GEN_14455;
      end
    end else begin
      cache_data_105 <= _GEN_14455;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h6a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_106 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_106 <= _GEN_14456;
      end
    end else begin
      cache_data_106 <= _GEN_14456;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h6b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_107 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_107 <= _GEN_14457;
      end
    end else begin
      cache_data_107 <= _GEN_14457;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h6c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_108 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_108 <= _GEN_14458;
      end
    end else begin
      cache_data_108 <= _GEN_14458;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h6d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_109 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_109 <= _GEN_14459;
      end
    end else begin
      cache_data_109 <= _GEN_14459;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h6e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_110 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_110 <= _GEN_14460;
      end
    end else begin
      cache_data_110 <= _GEN_14460;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h6f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_111 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_111 <= _GEN_14461;
      end
    end else begin
      cache_data_111 <= _GEN_14461;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h70 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_112 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_112 <= _GEN_14462;
      end
    end else begin
      cache_data_112 <= _GEN_14462;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h71 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_113 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_113 <= _GEN_14463;
      end
    end else begin
      cache_data_113 <= _GEN_14463;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h72 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_114 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_114 <= _GEN_14464;
      end
    end else begin
      cache_data_114 <= _GEN_14464;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h73 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_115 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_115 <= _GEN_14465;
      end
    end else begin
      cache_data_115 <= _GEN_14465;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h74 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_116 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_116 <= _GEN_14466;
      end
    end else begin
      cache_data_116 <= _GEN_14466;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h75 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_117 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_117 <= _GEN_14467;
      end
    end else begin
      cache_data_117 <= _GEN_14467;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h76 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_118 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_118 <= _GEN_14468;
      end
    end else begin
      cache_data_118 <= _GEN_14468;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h77 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_119 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_119 <= _GEN_14469;
      end
    end else begin
      cache_data_119 <= _GEN_14469;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h78 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_120 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_120 <= _GEN_14470;
      end
    end else begin
      cache_data_120 <= _GEN_14470;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h79 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_121 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_121 <= _GEN_14471;
      end
    end else begin
      cache_data_121 <= _GEN_14471;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h7a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_122 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_122 <= _GEN_14472;
      end
    end else begin
      cache_data_122 <= _GEN_14472;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h7b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_123 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_123 <= _GEN_14473;
      end
    end else begin
      cache_data_123 <= _GEN_14473;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h7c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_124 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_124 <= _GEN_14474;
      end
    end else begin
      cache_data_124 <= _GEN_14474;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h7d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_125 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_125 <= _GEN_14475;
      end
    end else begin
      cache_data_125 <= _GEN_14475;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h7e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_126 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_126 <= _GEN_14476;
      end
    end else begin
      cache_data_126 <= _GEN_14476;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h7f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_127 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_127 <= _GEN_14477;
      end
    end else begin
      cache_data_127 <= _GEN_14477;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h80 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_128 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_128 <= _GEN_14478;
      end
    end else begin
      cache_data_128 <= _GEN_14478;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h81 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_129 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_129 <= _GEN_14479;
      end
    end else begin
      cache_data_129 <= _GEN_14479;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h82 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_130 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_130 <= _GEN_14480;
      end
    end else begin
      cache_data_130 <= _GEN_14480;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h83 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_131 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_131 <= _GEN_14481;
      end
    end else begin
      cache_data_131 <= _GEN_14481;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h84 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_132 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_132 <= _GEN_14482;
      end
    end else begin
      cache_data_132 <= _GEN_14482;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h85 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_133 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_133 <= _GEN_14483;
      end
    end else begin
      cache_data_133 <= _GEN_14483;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h86 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_134 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_134 <= _GEN_14484;
      end
    end else begin
      cache_data_134 <= _GEN_14484;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h87 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_135 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_135 <= _GEN_14485;
      end
    end else begin
      cache_data_135 <= _GEN_14485;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h88 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_136 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_136 <= _GEN_14486;
      end
    end else begin
      cache_data_136 <= _GEN_14486;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h89 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_137 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_137 <= _GEN_14487;
      end
    end else begin
      cache_data_137 <= _GEN_14487;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h8a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_138 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_138 <= _GEN_14488;
      end
    end else begin
      cache_data_138 <= _GEN_14488;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h8b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_139 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_139 <= _GEN_14489;
      end
    end else begin
      cache_data_139 <= _GEN_14489;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h8c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_140 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_140 <= _GEN_14490;
      end
    end else begin
      cache_data_140 <= _GEN_14490;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h8d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_141 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_141 <= _GEN_14491;
      end
    end else begin
      cache_data_141 <= _GEN_14491;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h8e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_142 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_142 <= _GEN_14492;
      end
    end else begin
      cache_data_142 <= _GEN_14492;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h8f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_143 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_143 <= _GEN_14493;
      end
    end else begin
      cache_data_143 <= _GEN_14493;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h90 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_144 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_144 <= _GEN_14494;
      end
    end else begin
      cache_data_144 <= _GEN_14494;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h91 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_145 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_145 <= _GEN_14495;
      end
    end else begin
      cache_data_145 <= _GEN_14495;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h92 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_146 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_146 <= _GEN_14496;
      end
    end else begin
      cache_data_146 <= _GEN_14496;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h93 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_147 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_147 <= _GEN_14497;
      end
    end else begin
      cache_data_147 <= _GEN_14497;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h94 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_148 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_148 <= _GEN_14498;
      end
    end else begin
      cache_data_148 <= _GEN_14498;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h95 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_149 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_149 <= _GEN_14499;
      end
    end else begin
      cache_data_149 <= _GEN_14499;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h96 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_150 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_150 <= _GEN_14500;
      end
    end else begin
      cache_data_150 <= _GEN_14500;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h97 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_151 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_151 <= _GEN_14501;
      end
    end else begin
      cache_data_151 <= _GEN_14501;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h98 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_152 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_152 <= _GEN_14502;
      end
    end else begin
      cache_data_152 <= _GEN_14502;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h99 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_153 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_153 <= _GEN_14503;
      end
    end else begin
      cache_data_153 <= _GEN_14503;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h9a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_154 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_154 <= _GEN_14504;
      end
    end else begin
      cache_data_154 <= _GEN_14504;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h9b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_155 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_155 <= _GEN_14505;
      end
    end else begin
      cache_data_155 <= _GEN_14505;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h9c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_156 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_156 <= _GEN_14506;
      end
    end else begin
      cache_data_156 <= _GEN_14506;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h9d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_157 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_157 <= _GEN_14507;
      end
    end else begin
      cache_data_157 <= _GEN_14507;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h9e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_158 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_158 <= _GEN_14508;
      end
    end else begin
      cache_data_158 <= _GEN_14508;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h9f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_159 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_159 <= _GEN_14509;
      end
    end else begin
      cache_data_159 <= _GEN_14509;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'ha0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_160 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_160 <= _GEN_14510;
      end
    end else begin
      cache_data_160 <= _GEN_14510;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'ha1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_161 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_161 <= _GEN_14511;
      end
    end else begin
      cache_data_161 <= _GEN_14511;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'ha2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_162 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_162 <= _GEN_14512;
      end
    end else begin
      cache_data_162 <= _GEN_14512;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'ha3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_163 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_163 <= _GEN_14513;
      end
    end else begin
      cache_data_163 <= _GEN_14513;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'ha4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_164 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_164 <= _GEN_14514;
      end
    end else begin
      cache_data_164 <= _GEN_14514;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'ha5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_165 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_165 <= _GEN_14515;
      end
    end else begin
      cache_data_165 <= _GEN_14515;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'ha6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_166 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_166 <= _GEN_14516;
      end
    end else begin
      cache_data_166 <= _GEN_14516;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'ha7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_167 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_167 <= _GEN_14517;
      end
    end else begin
      cache_data_167 <= _GEN_14517;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'ha8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_168 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_168 <= _GEN_14518;
      end
    end else begin
      cache_data_168 <= _GEN_14518;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'ha9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_169 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_169 <= _GEN_14519;
      end
    end else begin
      cache_data_169 <= _GEN_14519;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'haa == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_170 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_170 <= _GEN_14520;
      end
    end else begin
      cache_data_170 <= _GEN_14520;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hab == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_171 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_171 <= _GEN_14521;
      end
    end else begin
      cache_data_171 <= _GEN_14521;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hac == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_172 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_172 <= _GEN_14522;
      end
    end else begin
      cache_data_172 <= _GEN_14522;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'had == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_173 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_173 <= _GEN_14523;
      end
    end else begin
      cache_data_173 <= _GEN_14523;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hae == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_174 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_174 <= _GEN_14524;
      end
    end else begin
      cache_data_174 <= _GEN_14524;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'haf == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_175 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_175 <= _GEN_14525;
      end
    end else begin
      cache_data_175 <= _GEN_14525;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hb0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_176 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_176 <= _GEN_14526;
      end
    end else begin
      cache_data_176 <= _GEN_14526;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hb1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_177 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_177 <= _GEN_14527;
      end
    end else begin
      cache_data_177 <= _GEN_14527;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hb2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_178 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_178 <= _GEN_14528;
      end
    end else begin
      cache_data_178 <= _GEN_14528;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hb3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_179 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_179 <= _GEN_14529;
      end
    end else begin
      cache_data_179 <= _GEN_14529;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hb4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_180 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_180 <= _GEN_14530;
      end
    end else begin
      cache_data_180 <= _GEN_14530;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hb5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_181 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_181 <= _GEN_14531;
      end
    end else begin
      cache_data_181 <= _GEN_14531;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hb6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_182 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_182 <= _GEN_14532;
      end
    end else begin
      cache_data_182 <= _GEN_14532;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hb7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_183 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_183 <= _GEN_14533;
      end
    end else begin
      cache_data_183 <= _GEN_14533;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hb8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_184 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_184 <= _GEN_14534;
      end
    end else begin
      cache_data_184 <= _GEN_14534;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hb9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_185 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_185 <= _GEN_14535;
      end
    end else begin
      cache_data_185 <= _GEN_14535;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hba == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_186 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_186 <= _GEN_14536;
      end
    end else begin
      cache_data_186 <= _GEN_14536;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hbb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_187 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_187 <= _GEN_14537;
      end
    end else begin
      cache_data_187 <= _GEN_14537;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hbc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_188 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_188 <= _GEN_14538;
      end
    end else begin
      cache_data_188 <= _GEN_14538;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hbd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_189 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_189 <= _GEN_14539;
      end
    end else begin
      cache_data_189 <= _GEN_14539;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hbe == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_190 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_190 <= _GEN_14540;
      end
    end else begin
      cache_data_190 <= _GEN_14540;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hbf == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_191 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_191 <= _GEN_14541;
      end
    end else begin
      cache_data_191 <= _GEN_14541;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hc0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_192 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_192 <= _GEN_14542;
      end
    end else begin
      cache_data_192 <= _GEN_14542;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hc1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_193 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_193 <= _GEN_14543;
      end
    end else begin
      cache_data_193 <= _GEN_14543;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hc2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_194 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_194 <= _GEN_14544;
      end
    end else begin
      cache_data_194 <= _GEN_14544;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hc3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_195 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_195 <= _GEN_14545;
      end
    end else begin
      cache_data_195 <= _GEN_14545;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hc4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_196 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_196 <= _GEN_14546;
      end
    end else begin
      cache_data_196 <= _GEN_14546;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hc5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_197 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_197 <= _GEN_14547;
      end
    end else begin
      cache_data_197 <= _GEN_14547;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hc6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_198 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_198 <= _GEN_14548;
      end
    end else begin
      cache_data_198 <= _GEN_14548;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hc7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_199 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_199 <= _GEN_14549;
      end
    end else begin
      cache_data_199 <= _GEN_14549;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hc8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_200 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_200 <= _GEN_14550;
      end
    end else begin
      cache_data_200 <= _GEN_14550;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hc9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_201 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_201 <= _GEN_14551;
      end
    end else begin
      cache_data_201 <= _GEN_14551;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hca == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_202 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_202 <= _GEN_14552;
      end
    end else begin
      cache_data_202 <= _GEN_14552;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hcb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_203 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_203 <= _GEN_14553;
      end
    end else begin
      cache_data_203 <= _GEN_14553;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hcc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_204 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_204 <= _GEN_14554;
      end
    end else begin
      cache_data_204 <= _GEN_14554;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hcd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_205 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_205 <= _GEN_14555;
      end
    end else begin
      cache_data_205 <= _GEN_14555;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hce == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_206 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_206 <= _GEN_14556;
      end
    end else begin
      cache_data_206 <= _GEN_14556;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hcf == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_207 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_207 <= _GEN_14557;
      end
    end else begin
      cache_data_207 <= _GEN_14557;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hd0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_208 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_208 <= _GEN_14558;
      end
    end else begin
      cache_data_208 <= _GEN_14558;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hd1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_209 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_209 <= _GEN_14559;
      end
    end else begin
      cache_data_209 <= _GEN_14559;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hd2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_210 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_210 <= _GEN_14560;
      end
    end else begin
      cache_data_210 <= _GEN_14560;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hd3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_211 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_211 <= _GEN_14561;
      end
    end else begin
      cache_data_211 <= _GEN_14561;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hd4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_212 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_212 <= _GEN_14562;
      end
    end else begin
      cache_data_212 <= _GEN_14562;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hd5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_213 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_213 <= _GEN_14563;
      end
    end else begin
      cache_data_213 <= _GEN_14563;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hd6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_214 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_214 <= _GEN_14564;
      end
    end else begin
      cache_data_214 <= _GEN_14564;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hd7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_215 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_215 <= _GEN_14565;
      end
    end else begin
      cache_data_215 <= _GEN_14565;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hd8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_216 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_216 <= _GEN_14566;
      end
    end else begin
      cache_data_216 <= _GEN_14566;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hd9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_217 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_217 <= _GEN_14567;
      end
    end else begin
      cache_data_217 <= _GEN_14567;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hda == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_218 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_218 <= _GEN_14568;
      end
    end else begin
      cache_data_218 <= _GEN_14568;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hdb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_219 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_219 <= _GEN_14569;
      end
    end else begin
      cache_data_219 <= _GEN_14569;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hdc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_220 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_220 <= _GEN_14570;
      end
    end else begin
      cache_data_220 <= _GEN_14570;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hdd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_221 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_221 <= _GEN_14571;
      end
    end else begin
      cache_data_221 <= _GEN_14571;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hde == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_222 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_222 <= _GEN_14572;
      end
    end else begin
      cache_data_222 <= _GEN_14572;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hdf == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_223 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_223 <= _GEN_14573;
      end
    end else begin
      cache_data_223 <= _GEN_14573;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'he0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_224 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_224 <= _GEN_14574;
      end
    end else begin
      cache_data_224 <= _GEN_14574;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'he1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_225 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_225 <= _GEN_14575;
      end
    end else begin
      cache_data_225 <= _GEN_14575;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'he2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_226 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_226 <= _GEN_14576;
      end
    end else begin
      cache_data_226 <= _GEN_14576;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'he3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_227 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_227 <= _GEN_14577;
      end
    end else begin
      cache_data_227 <= _GEN_14577;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'he4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_228 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_228 <= _GEN_14578;
      end
    end else begin
      cache_data_228 <= _GEN_14578;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'he5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_229 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_229 <= _GEN_14579;
      end
    end else begin
      cache_data_229 <= _GEN_14579;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'he6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_230 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_230 <= _GEN_14580;
      end
    end else begin
      cache_data_230 <= _GEN_14580;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'he7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_231 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_231 <= _GEN_14581;
      end
    end else begin
      cache_data_231 <= _GEN_14581;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'he8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_232 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_232 <= _GEN_14582;
      end
    end else begin
      cache_data_232 <= _GEN_14582;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'he9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_233 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_233 <= _GEN_14583;
      end
    end else begin
      cache_data_233 <= _GEN_14583;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hea == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_234 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_234 <= _GEN_14584;
      end
    end else begin
      cache_data_234 <= _GEN_14584;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'heb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_235 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_235 <= _GEN_14585;
      end
    end else begin
      cache_data_235 <= _GEN_14585;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hec == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_236 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_236 <= _GEN_14586;
      end
    end else begin
      cache_data_236 <= _GEN_14586;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hed == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_237 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_237 <= _GEN_14587;
      end
    end else begin
      cache_data_237 <= _GEN_14587;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hee == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_238 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_238 <= _GEN_14588;
      end
    end else begin
      cache_data_238 <= _GEN_14588;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hef == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_239 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_239 <= _GEN_14589;
      end
    end else begin
      cache_data_239 <= _GEN_14589;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hf0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_240 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_240 <= _GEN_14590;
      end
    end else begin
      cache_data_240 <= _GEN_14590;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hf1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_241 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_241 <= _GEN_14591;
      end
    end else begin
      cache_data_241 <= _GEN_14591;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hf2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_242 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_242 <= _GEN_14592;
      end
    end else begin
      cache_data_242 <= _GEN_14592;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hf3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_243 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_243 <= _GEN_14593;
      end
    end else begin
      cache_data_243 <= _GEN_14593;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hf4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_244 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_244 <= _GEN_14594;
      end
    end else begin
      cache_data_244 <= _GEN_14594;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hf5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_245 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_245 <= _GEN_14595;
      end
    end else begin
      cache_data_245 <= _GEN_14595;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hf6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_246 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_246 <= _GEN_14596;
      end
    end else begin
      cache_data_246 <= _GEN_14596;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hf7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_247 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_247 <= _GEN_14597;
      end
    end else begin
      cache_data_247 <= _GEN_14597;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hf8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_248 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_248 <= _GEN_14598;
      end
    end else begin
      cache_data_248 <= _GEN_14598;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hf9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_249 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_249 <= _GEN_14599;
      end
    end else begin
      cache_data_249 <= _GEN_14599;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hfa == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_250 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_250 <= _GEN_14600;
      end
    end else begin
      cache_data_250 <= _GEN_14600;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hfb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_251 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_251 <= _GEN_14601;
      end
    end else begin
      cache_data_251 <= _GEN_14601;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hfc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_252 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_252 <= _GEN_14602;
      end
    end else begin
      cache_data_252 <= _GEN_14602;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hfd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_253 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_253 <= _GEN_14603;
      end
    end else begin
      cache_data_253 <= _GEN_14603;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hfe == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_254 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_254 <= _GEN_14604;
      end
    end else begin
      cache_data_254 <= _GEN_14604;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'hff == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_255 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_255 <= _GEN_14605;
      end
    end else begin
      cache_data_255 <= _GEN_14605;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h100 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_256 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_256 <= _GEN_14606;
      end
    end else begin
      cache_data_256 <= _GEN_14606;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h101 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_257 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_257 <= _GEN_14607;
      end
    end else begin
      cache_data_257 <= _GEN_14607;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h102 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_258 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_258 <= _GEN_14608;
      end
    end else begin
      cache_data_258 <= _GEN_14608;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h103 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_259 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_259 <= _GEN_14609;
      end
    end else begin
      cache_data_259 <= _GEN_14609;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h104 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_260 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_260 <= _GEN_14610;
      end
    end else begin
      cache_data_260 <= _GEN_14610;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h105 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_261 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_261 <= _GEN_14611;
      end
    end else begin
      cache_data_261 <= _GEN_14611;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h106 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_262 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_262 <= _GEN_14612;
      end
    end else begin
      cache_data_262 <= _GEN_14612;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h107 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_263 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_263 <= _GEN_14613;
      end
    end else begin
      cache_data_263 <= _GEN_14613;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h108 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_264 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_264 <= _GEN_14614;
      end
    end else begin
      cache_data_264 <= _GEN_14614;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h109 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_265 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_265 <= _GEN_14615;
      end
    end else begin
      cache_data_265 <= _GEN_14615;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h10a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_266 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_266 <= _GEN_14616;
      end
    end else begin
      cache_data_266 <= _GEN_14616;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h10b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_267 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_267 <= _GEN_14617;
      end
    end else begin
      cache_data_267 <= _GEN_14617;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h10c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_268 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_268 <= _GEN_14618;
      end
    end else begin
      cache_data_268 <= _GEN_14618;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h10d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_269 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_269 <= _GEN_14619;
      end
    end else begin
      cache_data_269 <= _GEN_14619;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h10e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_270 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_270 <= _GEN_14620;
      end
    end else begin
      cache_data_270 <= _GEN_14620;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h10f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_271 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_271 <= _GEN_14621;
      end
    end else begin
      cache_data_271 <= _GEN_14621;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h110 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_272 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_272 <= _GEN_14622;
      end
    end else begin
      cache_data_272 <= _GEN_14622;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h111 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_273 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_273 <= _GEN_14623;
      end
    end else begin
      cache_data_273 <= _GEN_14623;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h112 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_274 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_274 <= _GEN_14624;
      end
    end else begin
      cache_data_274 <= _GEN_14624;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h113 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_275 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_275 <= _GEN_14625;
      end
    end else begin
      cache_data_275 <= _GEN_14625;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h114 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_276 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_276 <= _GEN_14626;
      end
    end else begin
      cache_data_276 <= _GEN_14626;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h115 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_277 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_277 <= _GEN_14627;
      end
    end else begin
      cache_data_277 <= _GEN_14627;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h116 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_278 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_278 <= _GEN_14628;
      end
    end else begin
      cache_data_278 <= _GEN_14628;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h117 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_279 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_279 <= _GEN_14629;
      end
    end else begin
      cache_data_279 <= _GEN_14629;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h118 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_280 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_280 <= _GEN_14630;
      end
    end else begin
      cache_data_280 <= _GEN_14630;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h119 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_281 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_281 <= _GEN_14631;
      end
    end else begin
      cache_data_281 <= _GEN_14631;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h11a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_282 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_282 <= _GEN_14632;
      end
    end else begin
      cache_data_282 <= _GEN_14632;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h11b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_283 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_283 <= _GEN_14633;
      end
    end else begin
      cache_data_283 <= _GEN_14633;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h11c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_284 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_284 <= _GEN_14634;
      end
    end else begin
      cache_data_284 <= _GEN_14634;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h11d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_285 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_285 <= _GEN_14635;
      end
    end else begin
      cache_data_285 <= _GEN_14635;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h11e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_286 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_286 <= _GEN_14636;
      end
    end else begin
      cache_data_286 <= _GEN_14636;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h11f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_287 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_287 <= _GEN_14637;
      end
    end else begin
      cache_data_287 <= _GEN_14637;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h120 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_288 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_288 <= _GEN_14638;
      end
    end else begin
      cache_data_288 <= _GEN_14638;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h121 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_289 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_289 <= _GEN_14639;
      end
    end else begin
      cache_data_289 <= _GEN_14639;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h122 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_290 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_290 <= _GEN_14640;
      end
    end else begin
      cache_data_290 <= _GEN_14640;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h123 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_291 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_291 <= _GEN_14641;
      end
    end else begin
      cache_data_291 <= _GEN_14641;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h124 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_292 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_292 <= _GEN_14642;
      end
    end else begin
      cache_data_292 <= _GEN_14642;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h125 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_293 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_293 <= _GEN_14643;
      end
    end else begin
      cache_data_293 <= _GEN_14643;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h126 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_294 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_294 <= _GEN_14644;
      end
    end else begin
      cache_data_294 <= _GEN_14644;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h127 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_295 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_295 <= _GEN_14645;
      end
    end else begin
      cache_data_295 <= _GEN_14645;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h128 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_296 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_296 <= _GEN_14646;
      end
    end else begin
      cache_data_296 <= _GEN_14646;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h129 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_297 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_297 <= _GEN_14647;
      end
    end else begin
      cache_data_297 <= _GEN_14647;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h12a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_298 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_298 <= _GEN_14648;
      end
    end else begin
      cache_data_298 <= _GEN_14648;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h12b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_299 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_299 <= _GEN_14649;
      end
    end else begin
      cache_data_299 <= _GEN_14649;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h12c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_300 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_300 <= _GEN_14650;
      end
    end else begin
      cache_data_300 <= _GEN_14650;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h12d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_301 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_301 <= _GEN_14651;
      end
    end else begin
      cache_data_301 <= _GEN_14651;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h12e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_302 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_302 <= _GEN_14652;
      end
    end else begin
      cache_data_302 <= _GEN_14652;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h12f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_303 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_303 <= _GEN_14653;
      end
    end else begin
      cache_data_303 <= _GEN_14653;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h130 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_304 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_304 <= _GEN_14654;
      end
    end else begin
      cache_data_304 <= _GEN_14654;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h131 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_305 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_305 <= _GEN_14655;
      end
    end else begin
      cache_data_305 <= _GEN_14655;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h132 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_306 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_306 <= _GEN_14656;
      end
    end else begin
      cache_data_306 <= _GEN_14656;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h133 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_307 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_307 <= _GEN_14657;
      end
    end else begin
      cache_data_307 <= _GEN_14657;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h134 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_308 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_308 <= _GEN_14658;
      end
    end else begin
      cache_data_308 <= _GEN_14658;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h135 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_309 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_309 <= _GEN_14659;
      end
    end else begin
      cache_data_309 <= _GEN_14659;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h136 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_310 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_310 <= _GEN_14660;
      end
    end else begin
      cache_data_310 <= _GEN_14660;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h137 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_311 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_311 <= _GEN_14661;
      end
    end else begin
      cache_data_311 <= _GEN_14661;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h138 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_312 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_312 <= _GEN_14662;
      end
    end else begin
      cache_data_312 <= _GEN_14662;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h139 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_313 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_313 <= _GEN_14663;
      end
    end else begin
      cache_data_313 <= _GEN_14663;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h13a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_314 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_314 <= _GEN_14664;
      end
    end else begin
      cache_data_314 <= _GEN_14664;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h13b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_315 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_315 <= _GEN_14665;
      end
    end else begin
      cache_data_315 <= _GEN_14665;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h13c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_316 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_316 <= _GEN_14666;
      end
    end else begin
      cache_data_316 <= _GEN_14666;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h13d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_317 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_317 <= _GEN_14667;
      end
    end else begin
      cache_data_317 <= _GEN_14667;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h13e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_318 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_318 <= _GEN_14668;
      end
    end else begin
      cache_data_318 <= _GEN_14668;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h13f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_319 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_319 <= _GEN_14669;
      end
    end else begin
      cache_data_319 <= _GEN_14669;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h140 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_320 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_320 <= _GEN_14670;
      end
    end else begin
      cache_data_320 <= _GEN_14670;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h141 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_321 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_321 <= _GEN_14671;
      end
    end else begin
      cache_data_321 <= _GEN_14671;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h142 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_322 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_322 <= _GEN_14672;
      end
    end else begin
      cache_data_322 <= _GEN_14672;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h143 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_323 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_323 <= _GEN_14673;
      end
    end else begin
      cache_data_323 <= _GEN_14673;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h144 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_324 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_324 <= _GEN_14674;
      end
    end else begin
      cache_data_324 <= _GEN_14674;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h145 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_325 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_325 <= _GEN_14675;
      end
    end else begin
      cache_data_325 <= _GEN_14675;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h146 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_326 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_326 <= _GEN_14676;
      end
    end else begin
      cache_data_326 <= _GEN_14676;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h147 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_327 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_327 <= _GEN_14677;
      end
    end else begin
      cache_data_327 <= _GEN_14677;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h148 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_328 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_328 <= _GEN_14678;
      end
    end else begin
      cache_data_328 <= _GEN_14678;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h149 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_329 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_329 <= _GEN_14679;
      end
    end else begin
      cache_data_329 <= _GEN_14679;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h14a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_330 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_330 <= _GEN_14680;
      end
    end else begin
      cache_data_330 <= _GEN_14680;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h14b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_331 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_331 <= _GEN_14681;
      end
    end else begin
      cache_data_331 <= _GEN_14681;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h14c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_332 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_332 <= _GEN_14682;
      end
    end else begin
      cache_data_332 <= _GEN_14682;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h14d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_333 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_333 <= _GEN_14683;
      end
    end else begin
      cache_data_333 <= _GEN_14683;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h14e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_334 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_334 <= _GEN_14684;
      end
    end else begin
      cache_data_334 <= _GEN_14684;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h14f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_335 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_335 <= _GEN_14685;
      end
    end else begin
      cache_data_335 <= _GEN_14685;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h150 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_336 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_336 <= _GEN_14686;
      end
    end else begin
      cache_data_336 <= _GEN_14686;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h151 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_337 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_337 <= _GEN_14687;
      end
    end else begin
      cache_data_337 <= _GEN_14687;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h152 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_338 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_338 <= _GEN_14688;
      end
    end else begin
      cache_data_338 <= _GEN_14688;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h153 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_339 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_339 <= _GEN_14689;
      end
    end else begin
      cache_data_339 <= _GEN_14689;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h154 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_340 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_340 <= _GEN_14690;
      end
    end else begin
      cache_data_340 <= _GEN_14690;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h155 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_341 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_341 <= _GEN_14691;
      end
    end else begin
      cache_data_341 <= _GEN_14691;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h156 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_342 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_342 <= _GEN_14692;
      end
    end else begin
      cache_data_342 <= _GEN_14692;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h157 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_343 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_343 <= _GEN_14693;
      end
    end else begin
      cache_data_343 <= _GEN_14693;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h158 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_344 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_344 <= _GEN_14694;
      end
    end else begin
      cache_data_344 <= _GEN_14694;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h159 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_345 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_345 <= _GEN_14695;
      end
    end else begin
      cache_data_345 <= _GEN_14695;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h15a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_346 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_346 <= _GEN_14696;
      end
    end else begin
      cache_data_346 <= _GEN_14696;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h15b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_347 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_347 <= _GEN_14697;
      end
    end else begin
      cache_data_347 <= _GEN_14697;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h15c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_348 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_348 <= _GEN_14698;
      end
    end else begin
      cache_data_348 <= _GEN_14698;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h15d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_349 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_349 <= _GEN_14699;
      end
    end else begin
      cache_data_349 <= _GEN_14699;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h15e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_350 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_350 <= _GEN_14700;
      end
    end else begin
      cache_data_350 <= _GEN_14700;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h15f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_351 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_351 <= _GEN_14701;
      end
    end else begin
      cache_data_351 <= _GEN_14701;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h160 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_352 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_352 <= _GEN_14702;
      end
    end else begin
      cache_data_352 <= _GEN_14702;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h161 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_353 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_353 <= _GEN_14703;
      end
    end else begin
      cache_data_353 <= _GEN_14703;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h162 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_354 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_354 <= _GEN_14704;
      end
    end else begin
      cache_data_354 <= _GEN_14704;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h163 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_355 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_355 <= _GEN_14705;
      end
    end else begin
      cache_data_355 <= _GEN_14705;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h164 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_356 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_356 <= _GEN_14706;
      end
    end else begin
      cache_data_356 <= _GEN_14706;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h165 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_357 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_357 <= _GEN_14707;
      end
    end else begin
      cache_data_357 <= _GEN_14707;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h166 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_358 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_358 <= _GEN_14708;
      end
    end else begin
      cache_data_358 <= _GEN_14708;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h167 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_359 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_359 <= _GEN_14709;
      end
    end else begin
      cache_data_359 <= _GEN_14709;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h168 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_360 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_360 <= _GEN_14710;
      end
    end else begin
      cache_data_360 <= _GEN_14710;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h169 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_361 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_361 <= _GEN_14711;
      end
    end else begin
      cache_data_361 <= _GEN_14711;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h16a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_362 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_362 <= _GEN_14712;
      end
    end else begin
      cache_data_362 <= _GEN_14712;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h16b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_363 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_363 <= _GEN_14713;
      end
    end else begin
      cache_data_363 <= _GEN_14713;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h16c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_364 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_364 <= _GEN_14714;
      end
    end else begin
      cache_data_364 <= _GEN_14714;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h16d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_365 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_365 <= _GEN_14715;
      end
    end else begin
      cache_data_365 <= _GEN_14715;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h16e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_366 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_366 <= _GEN_14716;
      end
    end else begin
      cache_data_366 <= _GEN_14716;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h16f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_367 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_367 <= _GEN_14717;
      end
    end else begin
      cache_data_367 <= _GEN_14717;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h170 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_368 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_368 <= _GEN_14718;
      end
    end else begin
      cache_data_368 <= _GEN_14718;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h171 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_369 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_369 <= _GEN_14719;
      end
    end else begin
      cache_data_369 <= _GEN_14719;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h172 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_370 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_370 <= _GEN_14720;
      end
    end else begin
      cache_data_370 <= _GEN_14720;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h173 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_371 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_371 <= _GEN_14721;
      end
    end else begin
      cache_data_371 <= _GEN_14721;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h174 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_372 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_372 <= _GEN_14722;
      end
    end else begin
      cache_data_372 <= _GEN_14722;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h175 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_373 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_373 <= _GEN_14723;
      end
    end else begin
      cache_data_373 <= _GEN_14723;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h176 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_374 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_374 <= _GEN_14724;
      end
    end else begin
      cache_data_374 <= _GEN_14724;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h177 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_375 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_375 <= _GEN_14725;
      end
    end else begin
      cache_data_375 <= _GEN_14725;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h178 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_376 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_376 <= _GEN_14726;
      end
    end else begin
      cache_data_376 <= _GEN_14726;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h179 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_377 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_377 <= _GEN_14727;
      end
    end else begin
      cache_data_377 <= _GEN_14727;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h17a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_378 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_378 <= _GEN_14728;
      end
    end else begin
      cache_data_378 <= _GEN_14728;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h17b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_379 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_379 <= _GEN_14729;
      end
    end else begin
      cache_data_379 <= _GEN_14729;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h17c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_380 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_380 <= _GEN_14730;
      end
    end else begin
      cache_data_380 <= _GEN_14730;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h17d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_381 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_381 <= _GEN_14731;
      end
    end else begin
      cache_data_381 <= _GEN_14731;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h17e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_382 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_382 <= _GEN_14732;
      end
    end else begin
      cache_data_382 <= _GEN_14732;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h17f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_383 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_383 <= _GEN_14733;
      end
    end else begin
      cache_data_383 <= _GEN_14733;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h180 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_384 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_384 <= _GEN_14734;
      end
    end else begin
      cache_data_384 <= _GEN_14734;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h181 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_385 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_385 <= _GEN_14735;
      end
    end else begin
      cache_data_385 <= _GEN_14735;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h182 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_386 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_386 <= _GEN_14736;
      end
    end else begin
      cache_data_386 <= _GEN_14736;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h183 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_387 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_387 <= _GEN_14737;
      end
    end else begin
      cache_data_387 <= _GEN_14737;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h184 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_388 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_388 <= _GEN_14738;
      end
    end else begin
      cache_data_388 <= _GEN_14738;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h185 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_389 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_389 <= _GEN_14739;
      end
    end else begin
      cache_data_389 <= _GEN_14739;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h186 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_390 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_390 <= _GEN_14740;
      end
    end else begin
      cache_data_390 <= _GEN_14740;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h187 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_391 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_391 <= _GEN_14741;
      end
    end else begin
      cache_data_391 <= _GEN_14741;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h188 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_392 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_392 <= _GEN_14742;
      end
    end else begin
      cache_data_392 <= _GEN_14742;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h189 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_393 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_393 <= _GEN_14743;
      end
    end else begin
      cache_data_393 <= _GEN_14743;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h18a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_394 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_394 <= _GEN_14744;
      end
    end else begin
      cache_data_394 <= _GEN_14744;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h18b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_395 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_395 <= _GEN_14745;
      end
    end else begin
      cache_data_395 <= _GEN_14745;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h18c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_396 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_396 <= _GEN_14746;
      end
    end else begin
      cache_data_396 <= _GEN_14746;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h18d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_397 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_397 <= _GEN_14747;
      end
    end else begin
      cache_data_397 <= _GEN_14747;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h18e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_398 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_398 <= _GEN_14748;
      end
    end else begin
      cache_data_398 <= _GEN_14748;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h18f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_399 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_399 <= _GEN_14749;
      end
    end else begin
      cache_data_399 <= _GEN_14749;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h190 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_400 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_400 <= _GEN_14750;
      end
    end else begin
      cache_data_400 <= _GEN_14750;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h191 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_401 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_401 <= _GEN_14751;
      end
    end else begin
      cache_data_401 <= _GEN_14751;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h192 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_402 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_402 <= _GEN_14752;
      end
    end else begin
      cache_data_402 <= _GEN_14752;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h193 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_403 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_403 <= _GEN_14753;
      end
    end else begin
      cache_data_403 <= _GEN_14753;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h194 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_404 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_404 <= _GEN_14754;
      end
    end else begin
      cache_data_404 <= _GEN_14754;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h195 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_405 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_405 <= _GEN_14755;
      end
    end else begin
      cache_data_405 <= _GEN_14755;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h196 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_406 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_406 <= _GEN_14756;
      end
    end else begin
      cache_data_406 <= _GEN_14756;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h197 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_407 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_407 <= _GEN_14757;
      end
    end else begin
      cache_data_407 <= _GEN_14757;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h198 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_408 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_408 <= _GEN_14758;
      end
    end else begin
      cache_data_408 <= _GEN_14758;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h199 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_409 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_409 <= _GEN_14759;
      end
    end else begin
      cache_data_409 <= _GEN_14759;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h19a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_410 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_410 <= _GEN_14760;
      end
    end else begin
      cache_data_410 <= _GEN_14760;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h19b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_411 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_411 <= _GEN_14761;
      end
    end else begin
      cache_data_411 <= _GEN_14761;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h19c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_412 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_412 <= _GEN_14762;
      end
    end else begin
      cache_data_412 <= _GEN_14762;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h19d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_413 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_413 <= _GEN_14763;
      end
    end else begin
      cache_data_413 <= _GEN_14763;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h19e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_414 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_414 <= _GEN_14764;
      end
    end else begin
      cache_data_414 <= _GEN_14764;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h19f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_415 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_415 <= _GEN_14765;
      end
    end else begin
      cache_data_415 <= _GEN_14765;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1a0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_416 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_416 <= _GEN_14766;
      end
    end else begin
      cache_data_416 <= _GEN_14766;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1a1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_417 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_417 <= _GEN_14767;
      end
    end else begin
      cache_data_417 <= _GEN_14767;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1a2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_418 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_418 <= _GEN_14768;
      end
    end else begin
      cache_data_418 <= _GEN_14768;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1a3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_419 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_419 <= _GEN_14769;
      end
    end else begin
      cache_data_419 <= _GEN_14769;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1a4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_420 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_420 <= _GEN_14770;
      end
    end else begin
      cache_data_420 <= _GEN_14770;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1a5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_421 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_421 <= _GEN_14771;
      end
    end else begin
      cache_data_421 <= _GEN_14771;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1a6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_422 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_422 <= _GEN_14772;
      end
    end else begin
      cache_data_422 <= _GEN_14772;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1a7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_423 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_423 <= _GEN_14773;
      end
    end else begin
      cache_data_423 <= _GEN_14773;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1a8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_424 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_424 <= _GEN_14774;
      end
    end else begin
      cache_data_424 <= _GEN_14774;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1a9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_425 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_425 <= _GEN_14775;
      end
    end else begin
      cache_data_425 <= _GEN_14775;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1aa == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_426 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_426 <= _GEN_14776;
      end
    end else begin
      cache_data_426 <= _GEN_14776;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ab == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_427 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_427 <= _GEN_14777;
      end
    end else begin
      cache_data_427 <= _GEN_14777;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ac == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_428 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_428 <= _GEN_14778;
      end
    end else begin
      cache_data_428 <= _GEN_14778;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ad == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_429 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_429 <= _GEN_14779;
      end
    end else begin
      cache_data_429 <= _GEN_14779;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ae == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_430 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_430 <= _GEN_14780;
      end
    end else begin
      cache_data_430 <= _GEN_14780;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1af == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_431 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_431 <= _GEN_14781;
      end
    end else begin
      cache_data_431 <= _GEN_14781;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1b0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_432 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_432 <= _GEN_14782;
      end
    end else begin
      cache_data_432 <= _GEN_14782;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1b1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_433 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_433 <= _GEN_14783;
      end
    end else begin
      cache_data_433 <= _GEN_14783;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1b2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_434 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_434 <= _GEN_14784;
      end
    end else begin
      cache_data_434 <= _GEN_14784;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1b3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_435 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_435 <= _GEN_14785;
      end
    end else begin
      cache_data_435 <= _GEN_14785;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1b4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_436 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_436 <= _GEN_14786;
      end
    end else begin
      cache_data_436 <= _GEN_14786;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1b5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_437 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_437 <= _GEN_14787;
      end
    end else begin
      cache_data_437 <= _GEN_14787;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1b6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_438 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_438 <= _GEN_14788;
      end
    end else begin
      cache_data_438 <= _GEN_14788;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1b7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_439 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_439 <= _GEN_14789;
      end
    end else begin
      cache_data_439 <= _GEN_14789;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1b8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_440 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_440 <= _GEN_14790;
      end
    end else begin
      cache_data_440 <= _GEN_14790;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1b9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_441 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_441 <= _GEN_14791;
      end
    end else begin
      cache_data_441 <= _GEN_14791;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ba == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_442 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_442 <= _GEN_14792;
      end
    end else begin
      cache_data_442 <= _GEN_14792;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1bb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_443 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_443 <= _GEN_14793;
      end
    end else begin
      cache_data_443 <= _GEN_14793;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1bc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_444 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_444 <= _GEN_14794;
      end
    end else begin
      cache_data_444 <= _GEN_14794;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1bd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_445 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_445 <= _GEN_14795;
      end
    end else begin
      cache_data_445 <= _GEN_14795;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1be == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_446 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_446 <= _GEN_14796;
      end
    end else begin
      cache_data_446 <= _GEN_14796;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1bf == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_447 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_447 <= _GEN_14797;
      end
    end else begin
      cache_data_447 <= _GEN_14797;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1c0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_448 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_448 <= _GEN_14798;
      end
    end else begin
      cache_data_448 <= _GEN_14798;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1c1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_449 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_449 <= _GEN_14799;
      end
    end else begin
      cache_data_449 <= _GEN_14799;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1c2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_450 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_450 <= _GEN_14800;
      end
    end else begin
      cache_data_450 <= _GEN_14800;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1c3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_451 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_451 <= _GEN_14801;
      end
    end else begin
      cache_data_451 <= _GEN_14801;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1c4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_452 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_452 <= _GEN_14802;
      end
    end else begin
      cache_data_452 <= _GEN_14802;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1c5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_453 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_453 <= _GEN_14803;
      end
    end else begin
      cache_data_453 <= _GEN_14803;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1c6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_454 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_454 <= _GEN_14804;
      end
    end else begin
      cache_data_454 <= _GEN_14804;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1c7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_455 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_455 <= _GEN_14805;
      end
    end else begin
      cache_data_455 <= _GEN_14805;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1c8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_456 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_456 <= _GEN_14806;
      end
    end else begin
      cache_data_456 <= _GEN_14806;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1c9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_457 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_457 <= _GEN_14807;
      end
    end else begin
      cache_data_457 <= _GEN_14807;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ca == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_458 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_458 <= _GEN_14808;
      end
    end else begin
      cache_data_458 <= _GEN_14808;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1cb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_459 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_459 <= _GEN_14809;
      end
    end else begin
      cache_data_459 <= _GEN_14809;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1cc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_460 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_460 <= _GEN_14810;
      end
    end else begin
      cache_data_460 <= _GEN_14810;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1cd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_461 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_461 <= _GEN_14811;
      end
    end else begin
      cache_data_461 <= _GEN_14811;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ce == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_462 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_462 <= _GEN_14812;
      end
    end else begin
      cache_data_462 <= _GEN_14812;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1cf == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_463 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_463 <= _GEN_14813;
      end
    end else begin
      cache_data_463 <= _GEN_14813;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1d0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_464 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_464 <= _GEN_14814;
      end
    end else begin
      cache_data_464 <= _GEN_14814;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1d1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_465 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_465 <= _GEN_14815;
      end
    end else begin
      cache_data_465 <= _GEN_14815;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1d2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_466 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_466 <= _GEN_14816;
      end
    end else begin
      cache_data_466 <= _GEN_14816;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1d3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_467 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_467 <= _GEN_14817;
      end
    end else begin
      cache_data_467 <= _GEN_14817;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1d4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_468 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_468 <= _GEN_14818;
      end
    end else begin
      cache_data_468 <= _GEN_14818;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1d5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_469 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_469 <= _GEN_14819;
      end
    end else begin
      cache_data_469 <= _GEN_14819;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1d6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_470 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_470 <= _GEN_14820;
      end
    end else begin
      cache_data_470 <= _GEN_14820;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1d7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_471 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_471 <= _GEN_14821;
      end
    end else begin
      cache_data_471 <= _GEN_14821;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1d8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_472 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_472 <= _GEN_14822;
      end
    end else begin
      cache_data_472 <= _GEN_14822;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1d9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_473 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_473 <= _GEN_14823;
      end
    end else begin
      cache_data_473 <= _GEN_14823;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1da == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_474 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_474 <= _GEN_14824;
      end
    end else begin
      cache_data_474 <= _GEN_14824;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1db == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_475 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_475 <= _GEN_14825;
      end
    end else begin
      cache_data_475 <= _GEN_14825;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1dc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_476 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_476 <= _GEN_14826;
      end
    end else begin
      cache_data_476 <= _GEN_14826;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1dd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_477 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_477 <= _GEN_14827;
      end
    end else begin
      cache_data_477 <= _GEN_14827;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1de == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_478 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_478 <= _GEN_14828;
      end
    end else begin
      cache_data_478 <= _GEN_14828;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1df == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_479 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_479 <= _GEN_14829;
      end
    end else begin
      cache_data_479 <= _GEN_14829;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1e0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_480 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_480 <= _GEN_14830;
      end
    end else begin
      cache_data_480 <= _GEN_14830;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1e1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_481 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_481 <= _GEN_14831;
      end
    end else begin
      cache_data_481 <= _GEN_14831;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1e2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_482 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_482 <= _GEN_14832;
      end
    end else begin
      cache_data_482 <= _GEN_14832;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1e3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_483 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_483 <= _GEN_14833;
      end
    end else begin
      cache_data_483 <= _GEN_14833;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1e4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_484 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_484 <= _GEN_14834;
      end
    end else begin
      cache_data_484 <= _GEN_14834;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1e5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_485 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_485 <= _GEN_14835;
      end
    end else begin
      cache_data_485 <= _GEN_14835;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1e6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_486 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_486 <= _GEN_14836;
      end
    end else begin
      cache_data_486 <= _GEN_14836;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1e7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_487 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_487 <= _GEN_14837;
      end
    end else begin
      cache_data_487 <= _GEN_14837;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1e8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_488 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_488 <= _GEN_14838;
      end
    end else begin
      cache_data_488 <= _GEN_14838;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1e9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_489 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_489 <= _GEN_14839;
      end
    end else begin
      cache_data_489 <= _GEN_14839;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ea == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_490 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_490 <= _GEN_14840;
      end
    end else begin
      cache_data_490 <= _GEN_14840;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1eb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_491 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_491 <= _GEN_14841;
      end
    end else begin
      cache_data_491 <= _GEN_14841;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ec == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_492 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_492 <= _GEN_14842;
      end
    end else begin
      cache_data_492 <= _GEN_14842;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ed == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_493 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_493 <= _GEN_14843;
      end
    end else begin
      cache_data_493 <= _GEN_14843;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ee == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_494 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_494 <= _GEN_14844;
      end
    end else begin
      cache_data_494 <= _GEN_14844;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ef == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_495 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_495 <= _GEN_14845;
      end
    end else begin
      cache_data_495 <= _GEN_14845;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1f0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_496 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_496 <= _GEN_14846;
      end
    end else begin
      cache_data_496 <= _GEN_14846;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1f1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_497 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_497 <= _GEN_14847;
      end
    end else begin
      cache_data_497 <= _GEN_14847;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1f2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_498 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_498 <= _GEN_14848;
      end
    end else begin
      cache_data_498 <= _GEN_14848;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1f3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_499 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_499 <= _GEN_14849;
      end
    end else begin
      cache_data_499 <= _GEN_14849;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1f4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_500 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_500 <= _GEN_14850;
      end
    end else begin
      cache_data_500 <= _GEN_14850;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1f5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_501 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_501 <= _GEN_14851;
      end
    end else begin
      cache_data_501 <= _GEN_14851;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1f6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_502 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_502 <= _GEN_14852;
      end
    end else begin
      cache_data_502 <= _GEN_14852;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1f7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_503 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_503 <= _GEN_14853;
      end
    end else begin
      cache_data_503 <= _GEN_14853;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1f8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_504 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_504 <= _GEN_14854;
      end
    end else begin
      cache_data_504 <= _GEN_14854;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1f9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_505 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_505 <= _GEN_14855;
      end
    end else begin
      cache_data_505 <= _GEN_14855;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1fa == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_506 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_506 <= _GEN_14856;
      end
    end else begin
      cache_data_506 <= _GEN_14856;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1fb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_507 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_507 <= _GEN_14857;
      end
    end else begin
      cache_data_507 <= _GEN_14857;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1fc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_508 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_508 <= _GEN_14858;
      end
    end else begin
      cache_data_508 <= _GEN_14858;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1fd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_509 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_509 <= _GEN_14859;
      end
    end else begin
      cache_data_509 <= _GEN_14859;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1fe == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_510 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_510 <= _GEN_14860;
      end
    end else begin
      cache_data_510 <= _GEN_14860;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h1ff == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_511 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_511 <= _GEN_14861;
      end
    end else begin
      cache_data_511 <= _GEN_14861;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h200 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_512 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_512 <= _GEN_14862;
      end
    end else begin
      cache_data_512 <= _GEN_14862;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h201 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_513 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_513 <= _GEN_14863;
      end
    end else begin
      cache_data_513 <= _GEN_14863;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h202 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_514 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_514 <= _GEN_14864;
      end
    end else begin
      cache_data_514 <= _GEN_14864;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h203 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_515 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_515 <= _GEN_14865;
      end
    end else begin
      cache_data_515 <= _GEN_14865;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h204 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_516 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_516 <= _GEN_14866;
      end
    end else begin
      cache_data_516 <= _GEN_14866;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h205 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_517 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_517 <= _GEN_14867;
      end
    end else begin
      cache_data_517 <= _GEN_14867;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h206 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_518 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_518 <= _GEN_14868;
      end
    end else begin
      cache_data_518 <= _GEN_14868;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h207 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_519 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_519 <= _GEN_14869;
      end
    end else begin
      cache_data_519 <= _GEN_14869;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h208 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_520 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_520 <= _GEN_14870;
      end
    end else begin
      cache_data_520 <= _GEN_14870;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h209 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_521 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_521 <= _GEN_14871;
      end
    end else begin
      cache_data_521 <= _GEN_14871;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h20a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_522 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_522 <= _GEN_14872;
      end
    end else begin
      cache_data_522 <= _GEN_14872;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h20b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_523 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_523 <= _GEN_14873;
      end
    end else begin
      cache_data_523 <= _GEN_14873;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h20c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_524 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_524 <= _GEN_14874;
      end
    end else begin
      cache_data_524 <= _GEN_14874;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h20d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_525 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_525 <= _GEN_14875;
      end
    end else begin
      cache_data_525 <= _GEN_14875;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h20e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_526 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_526 <= _GEN_14876;
      end
    end else begin
      cache_data_526 <= _GEN_14876;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h20f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_527 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_527 <= _GEN_14877;
      end
    end else begin
      cache_data_527 <= _GEN_14877;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h210 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_528 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_528 <= _GEN_14878;
      end
    end else begin
      cache_data_528 <= _GEN_14878;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h211 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_529 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_529 <= _GEN_14879;
      end
    end else begin
      cache_data_529 <= _GEN_14879;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h212 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_530 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_530 <= _GEN_14880;
      end
    end else begin
      cache_data_530 <= _GEN_14880;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h213 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_531 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_531 <= _GEN_14881;
      end
    end else begin
      cache_data_531 <= _GEN_14881;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h214 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_532 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_532 <= _GEN_14882;
      end
    end else begin
      cache_data_532 <= _GEN_14882;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h215 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_533 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_533 <= _GEN_14883;
      end
    end else begin
      cache_data_533 <= _GEN_14883;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h216 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_534 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_534 <= _GEN_14884;
      end
    end else begin
      cache_data_534 <= _GEN_14884;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h217 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_535 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_535 <= _GEN_14885;
      end
    end else begin
      cache_data_535 <= _GEN_14885;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h218 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_536 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_536 <= _GEN_14886;
      end
    end else begin
      cache_data_536 <= _GEN_14886;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h219 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_537 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_537 <= _GEN_14887;
      end
    end else begin
      cache_data_537 <= _GEN_14887;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h21a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_538 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_538 <= _GEN_14888;
      end
    end else begin
      cache_data_538 <= _GEN_14888;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h21b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_539 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_539 <= _GEN_14889;
      end
    end else begin
      cache_data_539 <= _GEN_14889;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h21c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_540 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_540 <= _GEN_14890;
      end
    end else begin
      cache_data_540 <= _GEN_14890;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h21d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_541 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_541 <= _GEN_14891;
      end
    end else begin
      cache_data_541 <= _GEN_14891;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h21e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_542 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_542 <= _GEN_14892;
      end
    end else begin
      cache_data_542 <= _GEN_14892;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h21f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_543 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_543 <= _GEN_14893;
      end
    end else begin
      cache_data_543 <= _GEN_14893;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h220 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_544 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_544 <= _GEN_14894;
      end
    end else begin
      cache_data_544 <= _GEN_14894;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h221 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_545 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_545 <= _GEN_14895;
      end
    end else begin
      cache_data_545 <= _GEN_14895;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h222 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_546 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_546 <= _GEN_14896;
      end
    end else begin
      cache_data_546 <= _GEN_14896;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h223 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_547 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_547 <= _GEN_14897;
      end
    end else begin
      cache_data_547 <= _GEN_14897;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h224 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_548 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_548 <= _GEN_14898;
      end
    end else begin
      cache_data_548 <= _GEN_14898;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h225 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_549 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_549 <= _GEN_14899;
      end
    end else begin
      cache_data_549 <= _GEN_14899;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h226 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_550 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_550 <= _GEN_14900;
      end
    end else begin
      cache_data_550 <= _GEN_14900;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h227 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_551 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_551 <= _GEN_14901;
      end
    end else begin
      cache_data_551 <= _GEN_14901;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h228 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_552 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_552 <= _GEN_14902;
      end
    end else begin
      cache_data_552 <= _GEN_14902;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h229 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_553 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_553 <= _GEN_14903;
      end
    end else begin
      cache_data_553 <= _GEN_14903;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h22a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_554 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_554 <= _GEN_14904;
      end
    end else begin
      cache_data_554 <= _GEN_14904;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h22b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_555 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_555 <= _GEN_14905;
      end
    end else begin
      cache_data_555 <= _GEN_14905;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h22c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_556 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_556 <= _GEN_14906;
      end
    end else begin
      cache_data_556 <= _GEN_14906;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h22d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_557 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_557 <= _GEN_14907;
      end
    end else begin
      cache_data_557 <= _GEN_14907;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h22e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_558 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_558 <= _GEN_14908;
      end
    end else begin
      cache_data_558 <= _GEN_14908;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h22f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_559 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_559 <= _GEN_14909;
      end
    end else begin
      cache_data_559 <= _GEN_14909;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h230 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_560 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_560 <= _GEN_14910;
      end
    end else begin
      cache_data_560 <= _GEN_14910;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h231 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_561 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_561 <= _GEN_14911;
      end
    end else begin
      cache_data_561 <= _GEN_14911;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h232 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_562 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_562 <= _GEN_14912;
      end
    end else begin
      cache_data_562 <= _GEN_14912;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h233 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_563 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_563 <= _GEN_14913;
      end
    end else begin
      cache_data_563 <= _GEN_14913;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h234 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_564 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_564 <= _GEN_14914;
      end
    end else begin
      cache_data_564 <= _GEN_14914;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h235 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_565 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_565 <= _GEN_14915;
      end
    end else begin
      cache_data_565 <= _GEN_14915;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h236 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_566 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_566 <= _GEN_14916;
      end
    end else begin
      cache_data_566 <= _GEN_14916;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h237 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_567 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_567 <= _GEN_14917;
      end
    end else begin
      cache_data_567 <= _GEN_14917;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h238 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_568 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_568 <= _GEN_14918;
      end
    end else begin
      cache_data_568 <= _GEN_14918;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h239 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_569 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_569 <= _GEN_14919;
      end
    end else begin
      cache_data_569 <= _GEN_14919;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h23a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_570 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_570 <= _GEN_14920;
      end
    end else begin
      cache_data_570 <= _GEN_14920;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h23b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_571 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_571 <= _GEN_14921;
      end
    end else begin
      cache_data_571 <= _GEN_14921;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h23c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_572 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_572 <= _GEN_14922;
      end
    end else begin
      cache_data_572 <= _GEN_14922;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h23d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_573 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_573 <= _GEN_14923;
      end
    end else begin
      cache_data_573 <= _GEN_14923;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h23e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_574 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_574 <= _GEN_14924;
      end
    end else begin
      cache_data_574 <= _GEN_14924;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h23f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_575 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_575 <= _GEN_14925;
      end
    end else begin
      cache_data_575 <= _GEN_14925;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h240 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_576 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_576 <= _GEN_14926;
      end
    end else begin
      cache_data_576 <= _GEN_14926;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h241 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_577 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_577 <= _GEN_14927;
      end
    end else begin
      cache_data_577 <= _GEN_14927;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h242 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_578 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_578 <= _GEN_14928;
      end
    end else begin
      cache_data_578 <= _GEN_14928;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h243 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_579 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_579 <= _GEN_14929;
      end
    end else begin
      cache_data_579 <= _GEN_14929;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h244 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_580 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_580 <= _GEN_14930;
      end
    end else begin
      cache_data_580 <= _GEN_14930;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h245 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_581 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_581 <= _GEN_14931;
      end
    end else begin
      cache_data_581 <= _GEN_14931;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h246 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_582 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_582 <= _GEN_14932;
      end
    end else begin
      cache_data_582 <= _GEN_14932;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h247 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_583 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_583 <= _GEN_14933;
      end
    end else begin
      cache_data_583 <= _GEN_14933;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h248 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_584 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_584 <= _GEN_14934;
      end
    end else begin
      cache_data_584 <= _GEN_14934;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h249 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_585 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_585 <= _GEN_14935;
      end
    end else begin
      cache_data_585 <= _GEN_14935;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h24a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_586 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_586 <= _GEN_14936;
      end
    end else begin
      cache_data_586 <= _GEN_14936;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h24b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_587 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_587 <= _GEN_14937;
      end
    end else begin
      cache_data_587 <= _GEN_14937;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h24c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_588 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_588 <= _GEN_14938;
      end
    end else begin
      cache_data_588 <= _GEN_14938;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h24d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_589 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_589 <= _GEN_14939;
      end
    end else begin
      cache_data_589 <= _GEN_14939;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h24e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_590 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_590 <= _GEN_14940;
      end
    end else begin
      cache_data_590 <= _GEN_14940;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h24f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_591 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_591 <= _GEN_14941;
      end
    end else begin
      cache_data_591 <= _GEN_14941;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h250 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_592 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_592 <= _GEN_14942;
      end
    end else begin
      cache_data_592 <= _GEN_14942;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h251 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_593 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_593 <= _GEN_14943;
      end
    end else begin
      cache_data_593 <= _GEN_14943;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h252 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_594 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_594 <= _GEN_14944;
      end
    end else begin
      cache_data_594 <= _GEN_14944;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h253 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_595 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_595 <= _GEN_14945;
      end
    end else begin
      cache_data_595 <= _GEN_14945;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h254 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_596 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_596 <= _GEN_14946;
      end
    end else begin
      cache_data_596 <= _GEN_14946;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h255 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_597 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_597 <= _GEN_14947;
      end
    end else begin
      cache_data_597 <= _GEN_14947;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h256 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_598 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_598 <= _GEN_14948;
      end
    end else begin
      cache_data_598 <= _GEN_14948;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h257 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_599 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_599 <= _GEN_14949;
      end
    end else begin
      cache_data_599 <= _GEN_14949;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h258 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_600 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_600 <= _GEN_14950;
      end
    end else begin
      cache_data_600 <= _GEN_14950;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h259 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_601 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_601 <= _GEN_14951;
      end
    end else begin
      cache_data_601 <= _GEN_14951;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h25a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_602 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_602 <= _GEN_14952;
      end
    end else begin
      cache_data_602 <= _GEN_14952;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h25b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_603 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_603 <= _GEN_14953;
      end
    end else begin
      cache_data_603 <= _GEN_14953;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h25c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_604 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_604 <= _GEN_14954;
      end
    end else begin
      cache_data_604 <= _GEN_14954;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h25d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_605 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_605 <= _GEN_14955;
      end
    end else begin
      cache_data_605 <= _GEN_14955;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h25e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_606 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_606 <= _GEN_14956;
      end
    end else begin
      cache_data_606 <= _GEN_14956;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h25f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_607 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_607 <= _GEN_14957;
      end
    end else begin
      cache_data_607 <= _GEN_14957;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h260 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_608 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_608 <= _GEN_14958;
      end
    end else begin
      cache_data_608 <= _GEN_14958;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h261 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_609 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_609 <= _GEN_14959;
      end
    end else begin
      cache_data_609 <= _GEN_14959;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h262 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_610 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_610 <= _GEN_14960;
      end
    end else begin
      cache_data_610 <= _GEN_14960;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h263 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_611 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_611 <= _GEN_14961;
      end
    end else begin
      cache_data_611 <= _GEN_14961;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h264 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_612 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_612 <= _GEN_14962;
      end
    end else begin
      cache_data_612 <= _GEN_14962;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h265 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_613 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_613 <= _GEN_14963;
      end
    end else begin
      cache_data_613 <= _GEN_14963;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h266 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_614 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_614 <= _GEN_14964;
      end
    end else begin
      cache_data_614 <= _GEN_14964;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h267 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_615 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_615 <= _GEN_14965;
      end
    end else begin
      cache_data_615 <= _GEN_14965;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h268 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_616 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_616 <= _GEN_14966;
      end
    end else begin
      cache_data_616 <= _GEN_14966;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h269 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_617 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_617 <= _GEN_14967;
      end
    end else begin
      cache_data_617 <= _GEN_14967;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h26a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_618 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_618 <= _GEN_14968;
      end
    end else begin
      cache_data_618 <= _GEN_14968;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h26b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_619 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_619 <= _GEN_14969;
      end
    end else begin
      cache_data_619 <= _GEN_14969;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h26c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_620 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_620 <= _GEN_14970;
      end
    end else begin
      cache_data_620 <= _GEN_14970;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h26d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_621 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_621 <= _GEN_14971;
      end
    end else begin
      cache_data_621 <= _GEN_14971;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h26e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_622 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_622 <= _GEN_14972;
      end
    end else begin
      cache_data_622 <= _GEN_14972;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h26f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_623 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_623 <= _GEN_14973;
      end
    end else begin
      cache_data_623 <= _GEN_14973;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h270 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_624 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_624 <= _GEN_14974;
      end
    end else begin
      cache_data_624 <= _GEN_14974;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h271 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_625 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_625 <= _GEN_14975;
      end
    end else begin
      cache_data_625 <= _GEN_14975;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h272 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_626 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_626 <= _GEN_14976;
      end
    end else begin
      cache_data_626 <= _GEN_14976;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h273 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_627 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_627 <= _GEN_14977;
      end
    end else begin
      cache_data_627 <= _GEN_14977;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h274 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_628 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_628 <= _GEN_14978;
      end
    end else begin
      cache_data_628 <= _GEN_14978;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h275 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_629 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_629 <= _GEN_14979;
      end
    end else begin
      cache_data_629 <= _GEN_14979;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h276 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_630 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_630 <= _GEN_14980;
      end
    end else begin
      cache_data_630 <= _GEN_14980;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h277 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_631 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_631 <= _GEN_14981;
      end
    end else begin
      cache_data_631 <= _GEN_14981;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h278 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_632 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_632 <= _GEN_14982;
      end
    end else begin
      cache_data_632 <= _GEN_14982;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h279 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_633 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_633 <= _GEN_14983;
      end
    end else begin
      cache_data_633 <= _GEN_14983;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h27a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_634 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_634 <= _GEN_14984;
      end
    end else begin
      cache_data_634 <= _GEN_14984;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h27b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_635 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_635 <= _GEN_14985;
      end
    end else begin
      cache_data_635 <= _GEN_14985;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h27c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_636 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_636 <= _GEN_14986;
      end
    end else begin
      cache_data_636 <= _GEN_14986;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h27d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_637 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_637 <= _GEN_14987;
      end
    end else begin
      cache_data_637 <= _GEN_14987;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h27e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_638 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_638 <= _GEN_14988;
      end
    end else begin
      cache_data_638 <= _GEN_14988;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h27f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_639 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_639 <= _GEN_14989;
      end
    end else begin
      cache_data_639 <= _GEN_14989;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h280 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_640 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_640 <= _GEN_14990;
      end
    end else begin
      cache_data_640 <= _GEN_14990;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h281 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_641 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_641 <= _GEN_14991;
      end
    end else begin
      cache_data_641 <= _GEN_14991;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h282 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_642 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_642 <= _GEN_14992;
      end
    end else begin
      cache_data_642 <= _GEN_14992;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h283 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_643 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_643 <= _GEN_14993;
      end
    end else begin
      cache_data_643 <= _GEN_14993;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h284 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_644 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_644 <= _GEN_14994;
      end
    end else begin
      cache_data_644 <= _GEN_14994;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h285 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_645 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_645 <= _GEN_14995;
      end
    end else begin
      cache_data_645 <= _GEN_14995;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h286 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_646 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_646 <= _GEN_14996;
      end
    end else begin
      cache_data_646 <= _GEN_14996;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h287 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_647 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_647 <= _GEN_14997;
      end
    end else begin
      cache_data_647 <= _GEN_14997;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h288 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_648 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_648 <= _GEN_14998;
      end
    end else begin
      cache_data_648 <= _GEN_14998;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h289 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_649 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_649 <= _GEN_14999;
      end
    end else begin
      cache_data_649 <= _GEN_14999;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h28a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_650 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_650 <= _GEN_15000;
      end
    end else begin
      cache_data_650 <= _GEN_15000;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h28b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_651 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_651 <= _GEN_15001;
      end
    end else begin
      cache_data_651 <= _GEN_15001;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h28c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_652 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_652 <= _GEN_15002;
      end
    end else begin
      cache_data_652 <= _GEN_15002;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h28d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_653 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_653 <= _GEN_15003;
      end
    end else begin
      cache_data_653 <= _GEN_15003;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h28e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_654 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_654 <= _GEN_15004;
      end
    end else begin
      cache_data_654 <= _GEN_15004;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h28f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_655 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_655 <= _GEN_15005;
      end
    end else begin
      cache_data_655 <= _GEN_15005;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h290 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_656 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_656 <= _GEN_15006;
      end
    end else begin
      cache_data_656 <= _GEN_15006;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h291 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_657 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_657 <= _GEN_15007;
      end
    end else begin
      cache_data_657 <= _GEN_15007;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h292 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_658 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_658 <= _GEN_15008;
      end
    end else begin
      cache_data_658 <= _GEN_15008;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h293 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_659 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_659 <= _GEN_15009;
      end
    end else begin
      cache_data_659 <= _GEN_15009;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h294 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_660 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_660 <= _GEN_15010;
      end
    end else begin
      cache_data_660 <= _GEN_15010;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h295 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_661 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_661 <= _GEN_15011;
      end
    end else begin
      cache_data_661 <= _GEN_15011;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h296 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_662 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_662 <= _GEN_15012;
      end
    end else begin
      cache_data_662 <= _GEN_15012;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h297 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_663 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_663 <= _GEN_15013;
      end
    end else begin
      cache_data_663 <= _GEN_15013;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h298 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_664 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_664 <= _GEN_15014;
      end
    end else begin
      cache_data_664 <= _GEN_15014;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h299 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_665 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_665 <= _GEN_15015;
      end
    end else begin
      cache_data_665 <= _GEN_15015;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h29a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_666 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_666 <= _GEN_15016;
      end
    end else begin
      cache_data_666 <= _GEN_15016;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h29b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_667 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_667 <= _GEN_15017;
      end
    end else begin
      cache_data_667 <= _GEN_15017;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h29c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_668 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_668 <= _GEN_15018;
      end
    end else begin
      cache_data_668 <= _GEN_15018;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h29d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_669 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_669 <= _GEN_15019;
      end
    end else begin
      cache_data_669 <= _GEN_15019;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h29e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_670 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_670 <= _GEN_15020;
      end
    end else begin
      cache_data_670 <= _GEN_15020;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h29f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_671 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_671 <= _GEN_15021;
      end
    end else begin
      cache_data_671 <= _GEN_15021;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2a0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_672 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_672 <= _GEN_15022;
      end
    end else begin
      cache_data_672 <= _GEN_15022;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2a1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_673 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_673 <= _GEN_15023;
      end
    end else begin
      cache_data_673 <= _GEN_15023;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2a2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_674 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_674 <= _GEN_15024;
      end
    end else begin
      cache_data_674 <= _GEN_15024;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2a3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_675 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_675 <= _GEN_15025;
      end
    end else begin
      cache_data_675 <= _GEN_15025;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2a4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_676 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_676 <= _GEN_15026;
      end
    end else begin
      cache_data_676 <= _GEN_15026;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2a5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_677 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_677 <= _GEN_15027;
      end
    end else begin
      cache_data_677 <= _GEN_15027;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2a6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_678 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_678 <= _GEN_15028;
      end
    end else begin
      cache_data_678 <= _GEN_15028;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2a7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_679 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_679 <= _GEN_15029;
      end
    end else begin
      cache_data_679 <= _GEN_15029;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2a8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_680 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_680 <= _GEN_15030;
      end
    end else begin
      cache_data_680 <= _GEN_15030;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2a9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_681 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_681 <= _GEN_15031;
      end
    end else begin
      cache_data_681 <= _GEN_15031;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2aa == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_682 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_682 <= _GEN_15032;
      end
    end else begin
      cache_data_682 <= _GEN_15032;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ab == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_683 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_683 <= _GEN_15033;
      end
    end else begin
      cache_data_683 <= _GEN_15033;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ac == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_684 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_684 <= _GEN_15034;
      end
    end else begin
      cache_data_684 <= _GEN_15034;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ad == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_685 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_685 <= _GEN_15035;
      end
    end else begin
      cache_data_685 <= _GEN_15035;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ae == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_686 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_686 <= _GEN_15036;
      end
    end else begin
      cache_data_686 <= _GEN_15036;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2af == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_687 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_687 <= _GEN_15037;
      end
    end else begin
      cache_data_687 <= _GEN_15037;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2b0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_688 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_688 <= _GEN_15038;
      end
    end else begin
      cache_data_688 <= _GEN_15038;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2b1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_689 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_689 <= _GEN_15039;
      end
    end else begin
      cache_data_689 <= _GEN_15039;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2b2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_690 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_690 <= _GEN_15040;
      end
    end else begin
      cache_data_690 <= _GEN_15040;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2b3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_691 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_691 <= _GEN_15041;
      end
    end else begin
      cache_data_691 <= _GEN_15041;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2b4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_692 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_692 <= _GEN_15042;
      end
    end else begin
      cache_data_692 <= _GEN_15042;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2b5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_693 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_693 <= _GEN_15043;
      end
    end else begin
      cache_data_693 <= _GEN_15043;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2b6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_694 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_694 <= _GEN_15044;
      end
    end else begin
      cache_data_694 <= _GEN_15044;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2b7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_695 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_695 <= _GEN_15045;
      end
    end else begin
      cache_data_695 <= _GEN_15045;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2b8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_696 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_696 <= _GEN_15046;
      end
    end else begin
      cache_data_696 <= _GEN_15046;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2b9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_697 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_697 <= _GEN_15047;
      end
    end else begin
      cache_data_697 <= _GEN_15047;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ba == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_698 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_698 <= _GEN_15048;
      end
    end else begin
      cache_data_698 <= _GEN_15048;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2bb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_699 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_699 <= _GEN_15049;
      end
    end else begin
      cache_data_699 <= _GEN_15049;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2bc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_700 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_700 <= _GEN_15050;
      end
    end else begin
      cache_data_700 <= _GEN_15050;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2bd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_701 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_701 <= _GEN_15051;
      end
    end else begin
      cache_data_701 <= _GEN_15051;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2be == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_702 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_702 <= _GEN_15052;
      end
    end else begin
      cache_data_702 <= _GEN_15052;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2bf == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_703 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_703 <= _GEN_15053;
      end
    end else begin
      cache_data_703 <= _GEN_15053;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2c0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_704 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_704 <= _GEN_15054;
      end
    end else begin
      cache_data_704 <= _GEN_15054;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2c1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_705 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_705 <= _GEN_15055;
      end
    end else begin
      cache_data_705 <= _GEN_15055;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2c2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_706 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_706 <= _GEN_15056;
      end
    end else begin
      cache_data_706 <= _GEN_15056;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2c3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_707 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_707 <= _GEN_15057;
      end
    end else begin
      cache_data_707 <= _GEN_15057;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2c4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_708 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_708 <= _GEN_15058;
      end
    end else begin
      cache_data_708 <= _GEN_15058;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2c5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_709 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_709 <= _GEN_15059;
      end
    end else begin
      cache_data_709 <= _GEN_15059;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2c6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_710 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_710 <= _GEN_15060;
      end
    end else begin
      cache_data_710 <= _GEN_15060;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2c7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_711 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_711 <= _GEN_15061;
      end
    end else begin
      cache_data_711 <= _GEN_15061;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2c8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_712 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_712 <= _GEN_15062;
      end
    end else begin
      cache_data_712 <= _GEN_15062;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2c9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_713 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_713 <= _GEN_15063;
      end
    end else begin
      cache_data_713 <= _GEN_15063;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ca == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_714 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_714 <= _GEN_15064;
      end
    end else begin
      cache_data_714 <= _GEN_15064;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2cb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_715 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_715 <= _GEN_15065;
      end
    end else begin
      cache_data_715 <= _GEN_15065;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2cc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_716 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_716 <= _GEN_15066;
      end
    end else begin
      cache_data_716 <= _GEN_15066;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2cd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_717 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_717 <= _GEN_15067;
      end
    end else begin
      cache_data_717 <= _GEN_15067;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ce == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_718 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_718 <= _GEN_15068;
      end
    end else begin
      cache_data_718 <= _GEN_15068;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2cf == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_719 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_719 <= _GEN_15069;
      end
    end else begin
      cache_data_719 <= _GEN_15069;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2d0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_720 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_720 <= _GEN_15070;
      end
    end else begin
      cache_data_720 <= _GEN_15070;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2d1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_721 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_721 <= _GEN_15071;
      end
    end else begin
      cache_data_721 <= _GEN_15071;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2d2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_722 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_722 <= _GEN_15072;
      end
    end else begin
      cache_data_722 <= _GEN_15072;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2d3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_723 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_723 <= _GEN_15073;
      end
    end else begin
      cache_data_723 <= _GEN_15073;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2d4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_724 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_724 <= _GEN_15074;
      end
    end else begin
      cache_data_724 <= _GEN_15074;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2d5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_725 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_725 <= _GEN_15075;
      end
    end else begin
      cache_data_725 <= _GEN_15075;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2d6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_726 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_726 <= _GEN_15076;
      end
    end else begin
      cache_data_726 <= _GEN_15076;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2d7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_727 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_727 <= _GEN_15077;
      end
    end else begin
      cache_data_727 <= _GEN_15077;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2d8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_728 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_728 <= _GEN_15078;
      end
    end else begin
      cache_data_728 <= _GEN_15078;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2d9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_729 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_729 <= _GEN_15079;
      end
    end else begin
      cache_data_729 <= _GEN_15079;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2da == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_730 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_730 <= _GEN_15080;
      end
    end else begin
      cache_data_730 <= _GEN_15080;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2db == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_731 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_731 <= _GEN_15081;
      end
    end else begin
      cache_data_731 <= _GEN_15081;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2dc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_732 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_732 <= _GEN_15082;
      end
    end else begin
      cache_data_732 <= _GEN_15082;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2dd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_733 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_733 <= _GEN_15083;
      end
    end else begin
      cache_data_733 <= _GEN_15083;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2de == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_734 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_734 <= _GEN_15084;
      end
    end else begin
      cache_data_734 <= _GEN_15084;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2df == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_735 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_735 <= _GEN_15085;
      end
    end else begin
      cache_data_735 <= _GEN_15085;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2e0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_736 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_736 <= _GEN_15086;
      end
    end else begin
      cache_data_736 <= _GEN_15086;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2e1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_737 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_737 <= _GEN_15087;
      end
    end else begin
      cache_data_737 <= _GEN_15087;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2e2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_738 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_738 <= _GEN_15088;
      end
    end else begin
      cache_data_738 <= _GEN_15088;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2e3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_739 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_739 <= _GEN_15089;
      end
    end else begin
      cache_data_739 <= _GEN_15089;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2e4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_740 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_740 <= _GEN_15090;
      end
    end else begin
      cache_data_740 <= _GEN_15090;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2e5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_741 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_741 <= _GEN_15091;
      end
    end else begin
      cache_data_741 <= _GEN_15091;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2e6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_742 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_742 <= _GEN_15092;
      end
    end else begin
      cache_data_742 <= _GEN_15092;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2e7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_743 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_743 <= _GEN_15093;
      end
    end else begin
      cache_data_743 <= _GEN_15093;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2e8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_744 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_744 <= _GEN_15094;
      end
    end else begin
      cache_data_744 <= _GEN_15094;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2e9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_745 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_745 <= _GEN_15095;
      end
    end else begin
      cache_data_745 <= _GEN_15095;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ea == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_746 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_746 <= _GEN_15096;
      end
    end else begin
      cache_data_746 <= _GEN_15096;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2eb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_747 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_747 <= _GEN_15097;
      end
    end else begin
      cache_data_747 <= _GEN_15097;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ec == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_748 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_748 <= _GEN_15098;
      end
    end else begin
      cache_data_748 <= _GEN_15098;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ed == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_749 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_749 <= _GEN_15099;
      end
    end else begin
      cache_data_749 <= _GEN_15099;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ee == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_750 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_750 <= _GEN_15100;
      end
    end else begin
      cache_data_750 <= _GEN_15100;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ef == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_751 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_751 <= _GEN_15101;
      end
    end else begin
      cache_data_751 <= _GEN_15101;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2f0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_752 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_752 <= _GEN_15102;
      end
    end else begin
      cache_data_752 <= _GEN_15102;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2f1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_753 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_753 <= _GEN_15103;
      end
    end else begin
      cache_data_753 <= _GEN_15103;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2f2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_754 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_754 <= _GEN_15104;
      end
    end else begin
      cache_data_754 <= _GEN_15104;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2f3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_755 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_755 <= _GEN_15105;
      end
    end else begin
      cache_data_755 <= _GEN_15105;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2f4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_756 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_756 <= _GEN_15106;
      end
    end else begin
      cache_data_756 <= _GEN_15106;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2f5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_757 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_757 <= _GEN_15107;
      end
    end else begin
      cache_data_757 <= _GEN_15107;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2f6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_758 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_758 <= _GEN_15108;
      end
    end else begin
      cache_data_758 <= _GEN_15108;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2f7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_759 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_759 <= _GEN_15109;
      end
    end else begin
      cache_data_759 <= _GEN_15109;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2f8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_760 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_760 <= _GEN_15110;
      end
    end else begin
      cache_data_760 <= _GEN_15110;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2f9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_761 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_761 <= _GEN_15111;
      end
    end else begin
      cache_data_761 <= _GEN_15111;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2fa == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_762 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_762 <= _GEN_15112;
      end
    end else begin
      cache_data_762 <= _GEN_15112;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2fb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_763 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_763 <= _GEN_15113;
      end
    end else begin
      cache_data_763 <= _GEN_15113;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2fc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_764 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_764 <= _GEN_15114;
      end
    end else begin
      cache_data_764 <= _GEN_15114;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2fd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_765 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_765 <= _GEN_15115;
      end
    end else begin
      cache_data_765 <= _GEN_15115;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2fe == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_766 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_766 <= _GEN_15116;
      end
    end else begin
      cache_data_766 <= _GEN_15116;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h2ff == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_767 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_767 <= _GEN_15117;
      end
    end else begin
      cache_data_767 <= _GEN_15117;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h300 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_768 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_768 <= _GEN_15118;
      end
    end else begin
      cache_data_768 <= _GEN_15118;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h301 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_769 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_769 <= _GEN_15119;
      end
    end else begin
      cache_data_769 <= _GEN_15119;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h302 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_770 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_770 <= _GEN_15120;
      end
    end else begin
      cache_data_770 <= _GEN_15120;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h303 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_771 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_771 <= _GEN_15121;
      end
    end else begin
      cache_data_771 <= _GEN_15121;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h304 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_772 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_772 <= _GEN_15122;
      end
    end else begin
      cache_data_772 <= _GEN_15122;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h305 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_773 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_773 <= _GEN_15123;
      end
    end else begin
      cache_data_773 <= _GEN_15123;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h306 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_774 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_774 <= _GEN_15124;
      end
    end else begin
      cache_data_774 <= _GEN_15124;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h307 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_775 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_775 <= _GEN_15125;
      end
    end else begin
      cache_data_775 <= _GEN_15125;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h308 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_776 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_776 <= _GEN_15126;
      end
    end else begin
      cache_data_776 <= _GEN_15126;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h309 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_777 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_777 <= _GEN_15127;
      end
    end else begin
      cache_data_777 <= _GEN_15127;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h30a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_778 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_778 <= _GEN_15128;
      end
    end else begin
      cache_data_778 <= _GEN_15128;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h30b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_779 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_779 <= _GEN_15129;
      end
    end else begin
      cache_data_779 <= _GEN_15129;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h30c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_780 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_780 <= _GEN_15130;
      end
    end else begin
      cache_data_780 <= _GEN_15130;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h30d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_781 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_781 <= _GEN_15131;
      end
    end else begin
      cache_data_781 <= _GEN_15131;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h30e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_782 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_782 <= _GEN_15132;
      end
    end else begin
      cache_data_782 <= _GEN_15132;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h30f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_783 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_783 <= _GEN_15133;
      end
    end else begin
      cache_data_783 <= _GEN_15133;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h310 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_784 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_784 <= _GEN_15134;
      end
    end else begin
      cache_data_784 <= _GEN_15134;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h311 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_785 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_785 <= _GEN_15135;
      end
    end else begin
      cache_data_785 <= _GEN_15135;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h312 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_786 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_786 <= _GEN_15136;
      end
    end else begin
      cache_data_786 <= _GEN_15136;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h313 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_787 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_787 <= _GEN_15137;
      end
    end else begin
      cache_data_787 <= _GEN_15137;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h314 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_788 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_788 <= _GEN_15138;
      end
    end else begin
      cache_data_788 <= _GEN_15138;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h315 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_789 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_789 <= _GEN_15139;
      end
    end else begin
      cache_data_789 <= _GEN_15139;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h316 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_790 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_790 <= _GEN_15140;
      end
    end else begin
      cache_data_790 <= _GEN_15140;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h317 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_791 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_791 <= _GEN_15141;
      end
    end else begin
      cache_data_791 <= _GEN_15141;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h318 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_792 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_792 <= _GEN_15142;
      end
    end else begin
      cache_data_792 <= _GEN_15142;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h319 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_793 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_793 <= _GEN_15143;
      end
    end else begin
      cache_data_793 <= _GEN_15143;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h31a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_794 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_794 <= _GEN_15144;
      end
    end else begin
      cache_data_794 <= _GEN_15144;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h31b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_795 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_795 <= _GEN_15145;
      end
    end else begin
      cache_data_795 <= _GEN_15145;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h31c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_796 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_796 <= _GEN_15146;
      end
    end else begin
      cache_data_796 <= _GEN_15146;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h31d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_797 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_797 <= _GEN_15147;
      end
    end else begin
      cache_data_797 <= _GEN_15147;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h31e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_798 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_798 <= _GEN_15148;
      end
    end else begin
      cache_data_798 <= _GEN_15148;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h31f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_799 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_799 <= _GEN_15149;
      end
    end else begin
      cache_data_799 <= _GEN_15149;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h320 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_800 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_800 <= _GEN_15150;
      end
    end else begin
      cache_data_800 <= _GEN_15150;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h321 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_801 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_801 <= _GEN_15151;
      end
    end else begin
      cache_data_801 <= _GEN_15151;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h322 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_802 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_802 <= _GEN_15152;
      end
    end else begin
      cache_data_802 <= _GEN_15152;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h323 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_803 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_803 <= _GEN_15153;
      end
    end else begin
      cache_data_803 <= _GEN_15153;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h324 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_804 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_804 <= _GEN_15154;
      end
    end else begin
      cache_data_804 <= _GEN_15154;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h325 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_805 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_805 <= _GEN_15155;
      end
    end else begin
      cache_data_805 <= _GEN_15155;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h326 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_806 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_806 <= _GEN_15156;
      end
    end else begin
      cache_data_806 <= _GEN_15156;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h327 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_807 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_807 <= _GEN_15157;
      end
    end else begin
      cache_data_807 <= _GEN_15157;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h328 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_808 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_808 <= _GEN_15158;
      end
    end else begin
      cache_data_808 <= _GEN_15158;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h329 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_809 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_809 <= _GEN_15159;
      end
    end else begin
      cache_data_809 <= _GEN_15159;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h32a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_810 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_810 <= _GEN_15160;
      end
    end else begin
      cache_data_810 <= _GEN_15160;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h32b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_811 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_811 <= _GEN_15161;
      end
    end else begin
      cache_data_811 <= _GEN_15161;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h32c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_812 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_812 <= _GEN_15162;
      end
    end else begin
      cache_data_812 <= _GEN_15162;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h32d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_813 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_813 <= _GEN_15163;
      end
    end else begin
      cache_data_813 <= _GEN_15163;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h32e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_814 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_814 <= _GEN_15164;
      end
    end else begin
      cache_data_814 <= _GEN_15164;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h32f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_815 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_815 <= _GEN_15165;
      end
    end else begin
      cache_data_815 <= _GEN_15165;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h330 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_816 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_816 <= _GEN_15166;
      end
    end else begin
      cache_data_816 <= _GEN_15166;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h331 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_817 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_817 <= _GEN_15167;
      end
    end else begin
      cache_data_817 <= _GEN_15167;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h332 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_818 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_818 <= _GEN_15168;
      end
    end else begin
      cache_data_818 <= _GEN_15168;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h333 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_819 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_819 <= _GEN_15169;
      end
    end else begin
      cache_data_819 <= _GEN_15169;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h334 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_820 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_820 <= _GEN_15170;
      end
    end else begin
      cache_data_820 <= _GEN_15170;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h335 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_821 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_821 <= _GEN_15171;
      end
    end else begin
      cache_data_821 <= _GEN_15171;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h336 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_822 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_822 <= _GEN_15172;
      end
    end else begin
      cache_data_822 <= _GEN_15172;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h337 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_823 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_823 <= _GEN_15173;
      end
    end else begin
      cache_data_823 <= _GEN_15173;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h338 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_824 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_824 <= _GEN_15174;
      end
    end else begin
      cache_data_824 <= _GEN_15174;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h339 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_825 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_825 <= _GEN_15175;
      end
    end else begin
      cache_data_825 <= _GEN_15175;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h33a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_826 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_826 <= _GEN_15176;
      end
    end else begin
      cache_data_826 <= _GEN_15176;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h33b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_827 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_827 <= _GEN_15177;
      end
    end else begin
      cache_data_827 <= _GEN_15177;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h33c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_828 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_828 <= _GEN_15178;
      end
    end else begin
      cache_data_828 <= _GEN_15178;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h33d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_829 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_829 <= _GEN_15179;
      end
    end else begin
      cache_data_829 <= _GEN_15179;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h33e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_830 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_830 <= _GEN_15180;
      end
    end else begin
      cache_data_830 <= _GEN_15180;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h33f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_831 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_831 <= _GEN_15181;
      end
    end else begin
      cache_data_831 <= _GEN_15181;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h340 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_832 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_832 <= _GEN_15182;
      end
    end else begin
      cache_data_832 <= _GEN_15182;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h341 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_833 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_833 <= _GEN_15183;
      end
    end else begin
      cache_data_833 <= _GEN_15183;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h342 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_834 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_834 <= _GEN_15184;
      end
    end else begin
      cache_data_834 <= _GEN_15184;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h343 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_835 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_835 <= _GEN_15185;
      end
    end else begin
      cache_data_835 <= _GEN_15185;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h344 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_836 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_836 <= _GEN_15186;
      end
    end else begin
      cache_data_836 <= _GEN_15186;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h345 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_837 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_837 <= _GEN_15187;
      end
    end else begin
      cache_data_837 <= _GEN_15187;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h346 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_838 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_838 <= _GEN_15188;
      end
    end else begin
      cache_data_838 <= _GEN_15188;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h347 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_839 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_839 <= _GEN_15189;
      end
    end else begin
      cache_data_839 <= _GEN_15189;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h348 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_840 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_840 <= _GEN_15190;
      end
    end else begin
      cache_data_840 <= _GEN_15190;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h349 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_841 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_841 <= _GEN_15191;
      end
    end else begin
      cache_data_841 <= _GEN_15191;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h34a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_842 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_842 <= _GEN_15192;
      end
    end else begin
      cache_data_842 <= _GEN_15192;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h34b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_843 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_843 <= _GEN_15193;
      end
    end else begin
      cache_data_843 <= _GEN_15193;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h34c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_844 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_844 <= _GEN_15194;
      end
    end else begin
      cache_data_844 <= _GEN_15194;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h34d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_845 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_845 <= _GEN_15195;
      end
    end else begin
      cache_data_845 <= _GEN_15195;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h34e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_846 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_846 <= _GEN_15196;
      end
    end else begin
      cache_data_846 <= _GEN_15196;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h34f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_847 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_847 <= _GEN_15197;
      end
    end else begin
      cache_data_847 <= _GEN_15197;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h350 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_848 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_848 <= _GEN_15198;
      end
    end else begin
      cache_data_848 <= _GEN_15198;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h351 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_849 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_849 <= _GEN_15199;
      end
    end else begin
      cache_data_849 <= _GEN_15199;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h352 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_850 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_850 <= _GEN_15200;
      end
    end else begin
      cache_data_850 <= _GEN_15200;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h353 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_851 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_851 <= _GEN_15201;
      end
    end else begin
      cache_data_851 <= _GEN_15201;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h354 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_852 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_852 <= _GEN_15202;
      end
    end else begin
      cache_data_852 <= _GEN_15202;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h355 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_853 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_853 <= _GEN_15203;
      end
    end else begin
      cache_data_853 <= _GEN_15203;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h356 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_854 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_854 <= _GEN_15204;
      end
    end else begin
      cache_data_854 <= _GEN_15204;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h357 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_855 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_855 <= _GEN_15205;
      end
    end else begin
      cache_data_855 <= _GEN_15205;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h358 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_856 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_856 <= _GEN_15206;
      end
    end else begin
      cache_data_856 <= _GEN_15206;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h359 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_857 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_857 <= _GEN_15207;
      end
    end else begin
      cache_data_857 <= _GEN_15207;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h35a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_858 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_858 <= _GEN_15208;
      end
    end else begin
      cache_data_858 <= _GEN_15208;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h35b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_859 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_859 <= _GEN_15209;
      end
    end else begin
      cache_data_859 <= _GEN_15209;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h35c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_860 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_860 <= _GEN_15210;
      end
    end else begin
      cache_data_860 <= _GEN_15210;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h35d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_861 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_861 <= _GEN_15211;
      end
    end else begin
      cache_data_861 <= _GEN_15211;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h35e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_862 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_862 <= _GEN_15212;
      end
    end else begin
      cache_data_862 <= _GEN_15212;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h35f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_863 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_863 <= _GEN_15213;
      end
    end else begin
      cache_data_863 <= _GEN_15213;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h360 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_864 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_864 <= _GEN_15214;
      end
    end else begin
      cache_data_864 <= _GEN_15214;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h361 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_865 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_865 <= _GEN_15215;
      end
    end else begin
      cache_data_865 <= _GEN_15215;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h362 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_866 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_866 <= _GEN_15216;
      end
    end else begin
      cache_data_866 <= _GEN_15216;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h363 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_867 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_867 <= _GEN_15217;
      end
    end else begin
      cache_data_867 <= _GEN_15217;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h364 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_868 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_868 <= _GEN_15218;
      end
    end else begin
      cache_data_868 <= _GEN_15218;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h365 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_869 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_869 <= _GEN_15219;
      end
    end else begin
      cache_data_869 <= _GEN_15219;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h366 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_870 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_870 <= _GEN_15220;
      end
    end else begin
      cache_data_870 <= _GEN_15220;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h367 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_871 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_871 <= _GEN_15221;
      end
    end else begin
      cache_data_871 <= _GEN_15221;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h368 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_872 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_872 <= _GEN_15222;
      end
    end else begin
      cache_data_872 <= _GEN_15222;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h369 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_873 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_873 <= _GEN_15223;
      end
    end else begin
      cache_data_873 <= _GEN_15223;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h36a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_874 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_874 <= _GEN_15224;
      end
    end else begin
      cache_data_874 <= _GEN_15224;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h36b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_875 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_875 <= _GEN_15225;
      end
    end else begin
      cache_data_875 <= _GEN_15225;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h36c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_876 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_876 <= _GEN_15226;
      end
    end else begin
      cache_data_876 <= _GEN_15226;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h36d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_877 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_877 <= _GEN_15227;
      end
    end else begin
      cache_data_877 <= _GEN_15227;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h36e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_878 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_878 <= _GEN_15228;
      end
    end else begin
      cache_data_878 <= _GEN_15228;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h36f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_879 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_879 <= _GEN_15229;
      end
    end else begin
      cache_data_879 <= _GEN_15229;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h370 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_880 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_880 <= _GEN_15230;
      end
    end else begin
      cache_data_880 <= _GEN_15230;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h371 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_881 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_881 <= _GEN_15231;
      end
    end else begin
      cache_data_881 <= _GEN_15231;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h372 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_882 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_882 <= _GEN_15232;
      end
    end else begin
      cache_data_882 <= _GEN_15232;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h373 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_883 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_883 <= _GEN_15233;
      end
    end else begin
      cache_data_883 <= _GEN_15233;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h374 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_884 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_884 <= _GEN_15234;
      end
    end else begin
      cache_data_884 <= _GEN_15234;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h375 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_885 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_885 <= _GEN_15235;
      end
    end else begin
      cache_data_885 <= _GEN_15235;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h376 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_886 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_886 <= _GEN_15236;
      end
    end else begin
      cache_data_886 <= _GEN_15236;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h377 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_887 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_887 <= _GEN_15237;
      end
    end else begin
      cache_data_887 <= _GEN_15237;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h378 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_888 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_888 <= _GEN_15238;
      end
    end else begin
      cache_data_888 <= _GEN_15238;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h379 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_889 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_889 <= _GEN_15239;
      end
    end else begin
      cache_data_889 <= _GEN_15239;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h37a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_890 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_890 <= _GEN_15240;
      end
    end else begin
      cache_data_890 <= _GEN_15240;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h37b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_891 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_891 <= _GEN_15241;
      end
    end else begin
      cache_data_891 <= _GEN_15241;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h37c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_892 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_892 <= _GEN_15242;
      end
    end else begin
      cache_data_892 <= _GEN_15242;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h37d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_893 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_893 <= _GEN_15243;
      end
    end else begin
      cache_data_893 <= _GEN_15243;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h37e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_894 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_894 <= _GEN_15244;
      end
    end else begin
      cache_data_894 <= _GEN_15244;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h37f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_895 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_895 <= _GEN_15245;
      end
    end else begin
      cache_data_895 <= _GEN_15245;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h380 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_896 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_896 <= _GEN_15246;
      end
    end else begin
      cache_data_896 <= _GEN_15246;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h381 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_897 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_897 <= _GEN_15247;
      end
    end else begin
      cache_data_897 <= _GEN_15247;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h382 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_898 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_898 <= _GEN_15248;
      end
    end else begin
      cache_data_898 <= _GEN_15248;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h383 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_899 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_899 <= _GEN_15249;
      end
    end else begin
      cache_data_899 <= _GEN_15249;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h384 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_900 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_900 <= _GEN_15250;
      end
    end else begin
      cache_data_900 <= _GEN_15250;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h385 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_901 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_901 <= _GEN_15251;
      end
    end else begin
      cache_data_901 <= _GEN_15251;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h386 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_902 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_902 <= _GEN_15252;
      end
    end else begin
      cache_data_902 <= _GEN_15252;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h387 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_903 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_903 <= _GEN_15253;
      end
    end else begin
      cache_data_903 <= _GEN_15253;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h388 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_904 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_904 <= _GEN_15254;
      end
    end else begin
      cache_data_904 <= _GEN_15254;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h389 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_905 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_905 <= _GEN_15255;
      end
    end else begin
      cache_data_905 <= _GEN_15255;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h38a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_906 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_906 <= _GEN_15256;
      end
    end else begin
      cache_data_906 <= _GEN_15256;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h38b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_907 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_907 <= _GEN_15257;
      end
    end else begin
      cache_data_907 <= _GEN_15257;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h38c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_908 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_908 <= _GEN_15258;
      end
    end else begin
      cache_data_908 <= _GEN_15258;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h38d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_909 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_909 <= _GEN_15259;
      end
    end else begin
      cache_data_909 <= _GEN_15259;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h38e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_910 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_910 <= _GEN_15260;
      end
    end else begin
      cache_data_910 <= _GEN_15260;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h38f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_911 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_911 <= _GEN_15261;
      end
    end else begin
      cache_data_911 <= _GEN_15261;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h390 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_912 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_912 <= _GEN_15262;
      end
    end else begin
      cache_data_912 <= _GEN_15262;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h391 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_913 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_913 <= _GEN_15263;
      end
    end else begin
      cache_data_913 <= _GEN_15263;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h392 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_914 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_914 <= _GEN_15264;
      end
    end else begin
      cache_data_914 <= _GEN_15264;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h393 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_915 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_915 <= _GEN_15265;
      end
    end else begin
      cache_data_915 <= _GEN_15265;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h394 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_916 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_916 <= _GEN_15266;
      end
    end else begin
      cache_data_916 <= _GEN_15266;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h395 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_917 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_917 <= _GEN_15267;
      end
    end else begin
      cache_data_917 <= _GEN_15267;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h396 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_918 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_918 <= _GEN_15268;
      end
    end else begin
      cache_data_918 <= _GEN_15268;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h397 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_919 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_919 <= _GEN_15269;
      end
    end else begin
      cache_data_919 <= _GEN_15269;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h398 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_920 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_920 <= _GEN_15270;
      end
    end else begin
      cache_data_920 <= _GEN_15270;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h399 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_921 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_921 <= _GEN_15271;
      end
    end else begin
      cache_data_921 <= _GEN_15271;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h39a == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_922 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_922 <= _GEN_15272;
      end
    end else begin
      cache_data_922 <= _GEN_15272;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h39b == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_923 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_923 <= _GEN_15273;
      end
    end else begin
      cache_data_923 <= _GEN_15273;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h39c == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_924 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_924 <= _GEN_15274;
      end
    end else begin
      cache_data_924 <= _GEN_15274;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h39d == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_925 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_925 <= _GEN_15275;
      end
    end else begin
      cache_data_925 <= _GEN_15275;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h39e == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_926 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_926 <= _GEN_15276;
      end
    end else begin
      cache_data_926 <= _GEN_15276;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h39f == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_927 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_927 <= _GEN_15277;
      end
    end else begin
      cache_data_927 <= _GEN_15277;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3a0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_928 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_928 <= _GEN_15278;
      end
    end else begin
      cache_data_928 <= _GEN_15278;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3a1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_929 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_929 <= _GEN_15279;
      end
    end else begin
      cache_data_929 <= _GEN_15279;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3a2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_930 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_930 <= _GEN_15280;
      end
    end else begin
      cache_data_930 <= _GEN_15280;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3a3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_931 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_931 <= _GEN_15281;
      end
    end else begin
      cache_data_931 <= _GEN_15281;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3a4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_932 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_932 <= _GEN_15282;
      end
    end else begin
      cache_data_932 <= _GEN_15282;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3a5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_933 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_933 <= _GEN_15283;
      end
    end else begin
      cache_data_933 <= _GEN_15283;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3a6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_934 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_934 <= _GEN_15284;
      end
    end else begin
      cache_data_934 <= _GEN_15284;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3a7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_935 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_935 <= _GEN_15285;
      end
    end else begin
      cache_data_935 <= _GEN_15285;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3a8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_936 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_936 <= _GEN_15286;
      end
    end else begin
      cache_data_936 <= _GEN_15286;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3a9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_937 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_937 <= _GEN_15287;
      end
    end else begin
      cache_data_937 <= _GEN_15287;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3aa == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_938 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_938 <= _GEN_15288;
      end
    end else begin
      cache_data_938 <= _GEN_15288;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ab == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_939 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_939 <= _GEN_15289;
      end
    end else begin
      cache_data_939 <= _GEN_15289;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ac == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_940 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_940 <= _GEN_15290;
      end
    end else begin
      cache_data_940 <= _GEN_15290;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ad == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_941 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_941 <= _GEN_15291;
      end
    end else begin
      cache_data_941 <= _GEN_15291;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ae == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_942 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_942 <= _GEN_15292;
      end
    end else begin
      cache_data_942 <= _GEN_15292;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3af == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_943 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_943 <= _GEN_15293;
      end
    end else begin
      cache_data_943 <= _GEN_15293;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3b0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_944 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_944 <= _GEN_15294;
      end
    end else begin
      cache_data_944 <= _GEN_15294;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3b1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_945 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_945 <= _GEN_15295;
      end
    end else begin
      cache_data_945 <= _GEN_15295;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3b2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_946 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_946 <= _GEN_15296;
      end
    end else begin
      cache_data_946 <= _GEN_15296;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3b3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_947 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_947 <= _GEN_15297;
      end
    end else begin
      cache_data_947 <= _GEN_15297;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3b4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_948 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_948 <= _GEN_15298;
      end
    end else begin
      cache_data_948 <= _GEN_15298;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3b5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_949 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_949 <= _GEN_15299;
      end
    end else begin
      cache_data_949 <= _GEN_15299;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3b6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_950 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_950 <= _GEN_15300;
      end
    end else begin
      cache_data_950 <= _GEN_15300;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3b7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_951 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_951 <= _GEN_15301;
      end
    end else begin
      cache_data_951 <= _GEN_15301;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3b8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_952 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_952 <= _GEN_15302;
      end
    end else begin
      cache_data_952 <= _GEN_15302;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3b9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_953 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_953 <= _GEN_15303;
      end
    end else begin
      cache_data_953 <= _GEN_15303;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ba == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_954 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_954 <= _GEN_15304;
      end
    end else begin
      cache_data_954 <= _GEN_15304;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3bb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_955 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_955 <= _GEN_15305;
      end
    end else begin
      cache_data_955 <= _GEN_15305;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3bc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_956 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_956 <= _GEN_15306;
      end
    end else begin
      cache_data_956 <= _GEN_15306;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3bd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_957 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_957 <= _GEN_15307;
      end
    end else begin
      cache_data_957 <= _GEN_15307;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3be == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_958 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_958 <= _GEN_15308;
      end
    end else begin
      cache_data_958 <= _GEN_15308;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3bf == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_959 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_959 <= _GEN_15309;
      end
    end else begin
      cache_data_959 <= _GEN_15309;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3c0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_960 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_960 <= _GEN_15310;
      end
    end else begin
      cache_data_960 <= _GEN_15310;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3c1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_961 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_961 <= _GEN_15311;
      end
    end else begin
      cache_data_961 <= _GEN_15311;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3c2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_962 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_962 <= _GEN_15312;
      end
    end else begin
      cache_data_962 <= _GEN_15312;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3c3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_963 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_963 <= _GEN_15313;
      end
    end else begin
      cache_data_963 <= _GEN_15313;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3c4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_964 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_964 <= _GEN_15314;
      end
    end else begin
      cache_data_964 <= _GEN_15314;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3c5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_965 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_965 <= _GEN_15315;
      end
    end else begin
      cache_data_965 <= _GEN_15315;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3c6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_966 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_966 <= _GEN_15316;
      end
    end else begin
      cache_data_966 <= _GEN_15316;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3c7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_967 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_967 <= _GEN_15317;
      end
    end else begin
      cache_data_967 <= _GEN_15317;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3c8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_968 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_968 <= _GEN_15318;
      end
    end else begin
      cache_data_968 <= _GEN_15318;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3c9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_969 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_969 <= _GEN_15319;
      end
    end else begin
      cache_data_969 <= _GEN_15319;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ca == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_970 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_970 <= _GEN_15320;
      end
    end else begin
      cache_data_970 <= _GEN_15320;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3cb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_971 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_971 <= _GEN_15321;
      end
    end else begin
      cache_data_971 <= _GEN_15321;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3cc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_972 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_972 <= _GEN_15322;
      end
    end else begin
      cache_data_972 <= _GEN_15322;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3cd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_973 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_973 <= _GEN_15323;
      end
    end else begin
      cache_data_973 <= _GEN_15323;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ce == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_974 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_974 <= _GEN_15324;
      end
    end else begin
      cache_data_974 <= _GEN_15324;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3cf == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_975 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_975 <= _GEN_15325;
      end
    end else begin
      cache_data_975 <= _GEN_15325;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3d0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_976 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_976 <= _GEN_15326;
      end
    end else begin
      cache_data_976 <= _GEN_15326;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3d1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_977 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_977 <= _GEN_15327;
      end
    end else begin
      cache_data_977 <= _GEN_15327;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3d2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_978 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_978 <= _GEN_15328;
      end
    end else begin
      cache_data_978 <= _GEN_15328;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3d3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_979 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_979 <= _GEN_15329;
      end
    end else begin
      cache_data_979 <= _GEN_15329;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3d4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_980 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_980 <= _GEN_15330;
      end
    end else begin
      cache_data_980 <= _GEN_15330;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3d5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_981 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_981 <= _GEN_15331;
      end
    end else begin
      cache_data_981 <= _GEN_15331;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3d6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_982 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_982 <= _GEN_15332;
      end
    end else begin
      cache_data_982 <= _GEN_15332;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3d7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_983 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_983 <= _GEN_15333;
      end
    end else begin
      cache_data_983 <= _GEN_15333;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3d8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_984 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_984 <= _GEN_15334;
      end
    end else begin
      cache_data_984 <= _GEN_15334;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3d9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_985 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_985 <= _GEN_15335;
      end
    end else begin
      cache_data_985 <= _GEN_15335;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3da == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_986 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_986 <= _GEN_15336;
      end
    end else begin
      cache_data_986 <= _GEN_15336;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3db == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_987 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_987 <= _GEN_15337;
      end
    end else begin
      cache_data_987 <= _GEN_15337;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3dc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_988 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_988 <= _GEN_15338;
      end
    end else begin
      cache_data_988 <= _GEN_15338;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3dd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_989 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_989 <= _GEN_15339;
      end
    end else begin
      cache_data_989 <= _GEN_15339;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3de == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_990 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_990 <= _GEN_15340;
      end
    end else begin
      cache_data_990 <= _GEN_15340;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3df == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_991 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_991 <= _GEN_15341;
      end
    end else begin
      cache_data_991 <= _GEN_15341;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3e0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_992 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_992 <= _GEN_15342;
      end
    end else begin
      cache_data_992 <= _GEN_15342;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3e1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_993 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_993 <= _GEN_15343;
      end
    end else begin
      cache_data_993 <= _GEN_15343;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3e2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_994 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_994 <= _GEN_15344;
      end
    end else begin
      cache_data_994 <= _GEN_15344;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3e3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_995 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_995 <= _GEN_15345;
      end
    end else begin
      cache_data_995 <= _GEN_15345;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3e4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_996 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_996 <= _GEN_15346;
      end
    end else begin
      cache_data_996 <= _GEN_15346;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3e5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_997 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_997 <= _GEN_15347;
      end
    end else begin
      cache_data_997 <= _GEN_15347;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3e6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_998 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_998 <= _GEN_15348;
      end
    end else begin
      cache_data_998 <= _GEN_15348;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3e7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_999 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_999 <= _GEN_15349;
      end
    end else begin
      cache_data_999 <= _GEN_15349;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3e8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1000 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1000 <= _GEN_15350;
      end
    end else begin
      cache_data_1000 <= _GEN_15350;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3e9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1001 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1001 <= _GEN_15351;
      end
    end else begin
      cache_data_1001 <= _GEN_15351;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ea == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1002 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1002 <= _GEN_15352;
      end
    end else begin
      cache_data_1002 <= _GEN_15352;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3eb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1003 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1003 <= _GEN_15353;
      end
    end else begin
      cache_data_1003 <= _GEN_15353;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ec == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1004 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1004 <= _GEN_15354;
      end
    end else begin
      cache_data_1004 <= _GEN_15354;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ed == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1005 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1005 <= _GEN_15355;
      end
    end else begin
      cache_data_1005 <= _GEN_15355;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ee == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1006 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1006 <= _GEN_15356;
      end
    end else begin
      cache_data_1006 <= _GEN_15356;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ef == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1007 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1007 <= _GEN_15357;
      end
    end else begin
      cache_data_1007 <= _GEN_15357;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3f0 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1008 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1008 <= _GEN_15358;
      end
    end else begin
      cache_data_1008 <= _GEN_15358;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3f1 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1009 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1009 <= _GEN_15359;
      end
    end else begin
      cache_data_1009 <= _GEN_15359;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3f2 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1010 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1010 <= _GEN_15360;
      end
    end else begin
      cache_data_1010 <= _GEN_15360;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3f3 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1011 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1011 <= _GEN_15361;
      end
    end else begin
      cache_data_1011 <= _GEN_15361;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3f4 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1012 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1012 <= _GEN_15362;
      end
    end else begin
      cache_data_1012 <= _GEN_15362;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3f5 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1013 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1013 <= _GEN_15363;
      end
    end else begin
      cache_data_1013 <= _GEN_15363;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3f6 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1014 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1014 <= _GEN_15364;
      end
    end else begin
      cache_data_1014 <= _GEN_15364;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3f7 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1015 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1015 <= _GEN_15365;
      end
    end else begin
      cache_data_1015 <= _GEN_15365;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3f8 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1016 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1016 <= _GEN_15366;
      end
    end else begin
      cache_data_1016 <= _GEN_15366;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3f9 == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1017 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1017 <= _GEN_15367;
      end
    end else begin
      cache_data_1017 <= _GEN_15367;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3fa == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1018 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1018 <= _GEN_15368;
      end
    end else begin
      cache_data_1018 <= _GEN_15368;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3fb == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1019 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1019 <= _GEN_15369;
      end
    end else begin
      cache_data_1019 <= _GEN_15369;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3fc == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1020 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1020 <= _GEN_15370;
      end
    end else begin
      cache_data_1020 <= _GEN_15370;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3fd == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1021 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1021 <= _GEN_15371;
      end
    end else begin
      cache_data_1021 <= _GEN_15371;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3fe == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1022 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1022 <= _GEN_15372;
      end
    end else begin
      cache_data_1022 <= _GEN_15372;
    end
    if (refill & io_inst_sram_data_ok) begin // @[icache.scala 141:41]
      if (10'h3ff == _dirty_T_1) begin // @[icache.scala 142:33]
        cache_data_1023 <= _cache_data_T_17; // @[icache.scala 142:33]
      end else begin
        cache_data_1023 <= _GEN_15373;
      end
    end else begin
      cache_data_1023 <= _GEN_15373;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  reg_rdata = _RAND_1[63:0];
  _RAND_2 = {1{`RANDOM}};
  delay = _RAND_2[0:0];
  _RAND_3 = {6{`RANDOM}};
  cache_data_0 = _RAND_3[184:0];
  _RAND_4 = {6{`RANDOM}};
  cache_data_1 = _RAND_4[184:0];
  _RAND_5 = {6{`RANDOM}};
  cache_data_2 = _RAND_5[184:0];
  _RAND_6 = {6{`RANDOM}};
  cache_data_3 = _RAND_6[184:0];
  _RAND_7 = {6{`RANDOM}};
  cache_data_4 = _RAND_7[184:0];
  _RAND_8 = {6{`RANDOM}};
  cache_data_5 = _RAND_8[184:0];
  _RAND_9 = {6{`RANDOM}};
  cache_data_6 = _RAND_9[184:0];
  _RAND_10 = {6{`RANDOM}};
  cache_data_7 = _RAND_10[184:0];
  _RAND_11 = {6{`RANDOM}};
  cache_data_8 = _RAND_11[184:0];
  _RAND_12 = {6{`RANDOM}};
  cache_data_9 = _RAND_12[184:0];
  _RAND_13 = {6{`RANDOM}};
  cache_data_10 = _RAND_13[184:0];
  _RAND_14 = {6{`RANDOM}};
  cache_data_11 = _RAND_14[184:0];
  _RAND_15 = {6{`RANDOM}};
  cache_data_12 = _RAND_15[184:0];
  _RAND_16 = {6{`RANDOM}};
  cache_data_13 = _RAND_16[184:0];
  _RAND_17 = {6{`RANDOM}};
  cache_data_14 = _RAND_17[184:0];
  _RAND_18 = {6{`RANDOM}};
  cache_data_15 = _RAND_18[184:0];
  _RAND_19 = {6{`RANDOM}};
  cache_data_16 = _RAND_19[184:0];
  _RAND_20 = {6{`RANDOM}};
  cache_data_17 = _RAND_20[184:0];
  _RAND_21 = {6{`RANDOM}};
  cache_data_18 = _RAND_21[184:0];
  _RAND_22 = {6{`RANDOM}};
  cache_data_19 = _RAND_22[184:0];
  _RAND_23 = {6{`RANDOM}};
  cache_data_20 = _RAND_23[184:0];
  _RAND_24 = {6{`RANDOM}};
  cache_data_21 = _RAND_24[184:0];
  _RAND_25 = {6{`RANDOM}};
  cache_data_22 = _RAND_25[184:0];
  _RAND_26 = {6{`RANDOM}};
  cache_data_23 = _RAND_26[184:0];
  _RAND_27 = {6{`RANDOM}};
  cache_data_24 = _RAND_27[184:0];
  _RAND_28 = {6{`RANDOM}};
  cache_data_25 = _RAND_28[184:0];
  _RAND_29 = {6{`RANDOM}};
  cache_data_26 = _RAND_29[184:0];
  _RAND_30 = {6{`RANDOM}};
  cache_data_27 = _RAND_30[184:0];
  _RAND_31 = {6{`RANDOM}};
  cache_data_28 = _RAND_31[184:0];
  _RAND_32 = {6{`RANDOM}};
  cache_data_29 = _RAND_32[184:0];
  _RAND_33 = {6{`RANDOM}};
  cache_data_30 = _RAND_33[184:0];
  _RAND_34 = {6{`RANDOM}};
  cache_data_31 = _RAND_34[184:0];
  _RAND_35 = {6{`RANDOM}};
  cache_data_32 = _RAND_35[184:0];
  _RAND_36 = {6{`RANDOM}};
  cache_data_33 = _RAND_36[184:0];
  _RAND_37 = {6{`RANDOM}};
  cache_data_34 = _RAND_37[184:0];
  _RAND_38 = {6{`RANDOM}};
  cache_data_35 = _RAND_38[184:0];
  _RAND_39 = {6{`RANDOM}};
  cache_data_36 = _RAND_39[184:0];
  _RAND_40 = {6{`RANDOM}};
  cache_data_37 = _RAND_40[184:0];
  _RAND_41 = {6{`RANDOM}};
  cache_data_38 = _RAND_41[184:0];
  _RAND_42 = {6{`RANDOM}};
  cache_data_39 = _RAND_42[184:0];
  _RAND_43 = {6{`RANDOM}};
  cache_data_40 = _RAND_43[184:0];
  _RAND_44 = {6{`RANDOM}};
  cache_data_41 = _RAND_44[184:0];
  _RAND_45 = {6{`RANDOM}};
  cache_data_42 = _RAND_45[184:0];
  _RAND_46 = {6{`RANDOM}};
  cache_data_43 = _RAND_46[184:0];
  _RAND_47 = {6{`RANDOM}};
  cache_data_44 = _RAND_47[184:0];
  _RAND_48 = {6{`RANDOM}};
  cache_data_45 = _RAND_48[184:0];
  _RAND_49 = {6{`RANDOM}};
  cache_data_46 = _RAND_49[184:0];
  _RAND_50 = {6{`RANDOM}};
  cache_data_47 = _RAND_50[184:0];
  _RAND_51 = {6{`RANDOM}};
  cache_data_48 = _RAND_51[184:0];
  _RAND_52 = {6{`RANDOM}};
  cache_data_49 = _RAND_52[184:0];
  _RAND_53 = {6{`RANDOM}};
  cache_data_50 = _RAND_53[184:0];
  _RAND_54 = {6{`RANDOM}};
  cache_data_51 = _RAND_54[184:0];
  _RAND_55 = {6{`RANDOM}};
  cache_data_52 = _RAND_55[184:0];
  _RAND_56 = {6{`RANDOM}};
  cache_data_53 = _RAND_56[184:0];
  _RAND_57 = {6{`RANDOM}};
  cache_data_54 = _RAND_57[184:0];
  _RAND_58 = {6{`RANDOM}};
  cache_data_55 = _RAND_58[184:0];
  _RAND_59 = {6{`RANDOM}};
  cache_data_56 = _RAND_59[184:0];
  _RAND_60 = {6{`RANDOM}};
  cache_data_57 = _RAND_60[184:0];
  _RAND_61 = {6{`RANDOM}};
  cache_data_58 = _RAND_61[184:0];
  _RAND_62 = {6{`RANDOM}};
  cache_data_59 = _RAND_62[184:0];
  _RAND_63 = {6{`RANDOM}};
  cache_data_60 = _RAND_63[184:0];
  _RAND_64 = {6{`RANDOM}};
  cache_data_61 = _RAND_64[184:0];
  _RAND_65 = {6{`RANDOM}};
  cache_data_62 = _RAND_65[184:0];
  _RAND_66 = {6{`RANDOM}};
  cache_data_63 = _RAND_66[184:0];
  _RAND_67 = {6{`RANDOM}};
  cache_data_64 = _RAND_67[184:0];
  _RAND_68 = {6{`RANDOM}};
  cache_data_65 = _RAND_68[184:0];
  _RAND_69 = {6{`RANDOM}};
  cache_data_66 = _RAND_69[184:0];
  _RAND_70 = {6{`RANDOM}};
  cache_data_67 = _RAND_70[184:0];
  _RAND_71 = {6{`RANDOM}};
  cache_data_68 = _RAND_71[184:0];
  _RAND_72 = {6{`RANDOM}};
  cache_data_69 = _RAND_72[184:0];
  _RAND_73 = {6{`RANDOM}};
  cache_data_70 = _RAND_73[184:0];
  _RAND_74 = {6{`RANDOM}};
  cache_data_71 = _RAND_74[184:0];
  _RAND_75 = {6{`RANDOM}};
  cache_data_72 = _RAND_75[184:0];
  _RAND_76 = {6{`RANDOM}};
  cache_data_73 = _RAND_76[184:0];
  _RAND_77 = {6{`RANDOM}};
  cache_data_74 = _RAND_77[184:0];
  _RAND_78 = {6{`RANDOM}};
  cache_data_75 = _RAND_78[184:0];
  _RAND_79 = {6{`RANDOM}};
  cache_data_76 = _RAND_79[184:0];
  _RAND_80 = {6{`RANDOM}};
  cache_data_77 = _RAND_80[184:0];
  _RAND_81 = {6{`RANDOM}};
  cache_data_78 = _RAND_81[184:0];
  _RAND_82 = {6{`RANDOM}};
  cache_data_79 = _RAND_82[184:0];
  _RAND_83 = {6{`RANDOM}};
  cache_data_80 = _RAND_83[184:0];
  _RAND_84 = {6{`RANDOM}};
  cache_data_81 = _RAND_84[184:0];
  _RAND_85 = {6{`RANDOM}};
  cache_data_82 = _RAND_85[184:0];
  _RAND_86 = {6{`RANDOM}};
  cache_data_83 = _RAND_86[184:0];
  _RAND_87 = {6{`RANDOM}};
  cache_data_84 = _RAND_87[184:0];
  _RAND_88 = {6{`RANDOM}};
  cache_data_85 = _RAND_88[184:0];
  _RAND_89 = {6{`RANDOM}};
  cache_data_86 = _RAND_89[184:0];
  _RAND_90 = {6{`RANDOM}};
  cache_data_87 = _RAND_90[184:0];
  _RAND_91 = {6{`RANDOM}};
  cache_data_88 = _RAND_91[184:0];
  _RAND_92 = {6{`RANDOM}};
  cache_data_89 = _RAND_92[184:0];
  _RAND_93 = {6{`RANDOM}};
  cache_data_90 = _RAND_93[184:0];
  _RAND_94 = {6{`RANDOM}};
  cache_data_91 = _RAND_94[184:0];
  _RAND_95 = {6{`RANDOM}};
  cache_data_92 = _RAND_95[184:0];
  _RAND_96 = {6{`RANDOM}};
  cache_data_93 = _RAND_96[184:0];
  _RAND_97 = {6{`RANDOM}};
  cache_data_94 = _RAND_97[184:0];
  _RAND_98 = {6{`RANDOM}};
  cache_data_95 = _RAND_98[184:0];
  _RAND_99 = {6{`RANDOM}};
  cache_data_96 = _RAND_99[184:0];
  _RAND_100 = {6{`RANDOM}};
  cache_data_97 = _RAND_100[184:0];
  _RAND_101 = {6{`RANDOM}};
  cache_data_98 = _RAND_101[184:0];
  _RAND_102 = {6{`RANDOM}};
  cache_data_99 = _RAND_102[184:0];
  _RAND_103 = {6{`RANDOM}};
  cache_data_100 = _RAND_103[184:0];
  _RAND_104 = {6{`RANDOM}};
  cache_data_101 = _RAND_104[184:0];
  _RAND_105 = {6{`RANDOM}};
  cache_data_102 = _RAND_105[184:0];
  _RAND_106 = {6{`RANDOM}};
  cache_data_103 = _RAND_106[184:0];
  _RAND_107 = {6{`RANDOM}};
  cache_data_104 = _RAND_107[184:0];
  _RAND_108 = {6{`RANDOM}};
  cache_data_105 = _RAND_108[184:0];
  _RAND_109 = {6{`RANDOM}};
  cache_data_106 = _RAND_109[184:0];
  _RAND_110 = {6{`RANDOM}};
  cache_data_107 = _RAND_110[184:0];
  _RAND_111 = {6{`RANDOM}};
  cache_data_108 = _RAND_111[184:0];
  _RAND_112 = {6{`RANDOM}};
  cache_data_109 = _RAND_112[184:0];
  _RAND_113 = {6{`RANDOM}};
  cache_data_110 = _RAND_113[184:0];
  _RAND_114 = {6{`RANDOM}};
  cache_data_111 = _RAND_114[184:0];
  _RAND_115 = {6{`RANDOM}};
  cache_data_112 = _RAND_115[184:0];
  _RAND_116 = {6{`RANDOM}};
  cache_data_113 = _RAND_116[184:0];
  _RAND_117 = {6{`RANDOM}};
  cache_data_114 = _RAND_117[184:0];
  _RAND_118 = {6{`RANDOM}};
  cache_data_115 = _RAND_118[184:0];
  _RAND_119 = {6{`RANDOM}};
  cache_data_116 = _RAND_119[184:0];
  _RAND_120 = {6{`RANDOM}};
  cache_data_117 = _RAND_120[184:0];
  _RAND_121 = {6{`RANDOM}};
  cache_data_118 = _RAND_121[184:0];
  _RAND_122 = {6{`RANDOM}};
  cache_data_119 = _RAND_122[184:0];
  _RAND_123 = {6{`RANDOM}};
  cache_data_120 = _RAND_123[184:0];
  _RAND_124 = {6{`RANDOM}};
  cache_data_121 = _RAND_124[184:0];
  _RAND_125 = {6{`RANDOM}};
  cache_data_122 = _RAND_125[184:0];
  _RAND_126 = {6{`RANDOM}};
  cache_data_123 = _RAND_126[184:0];
  _RAND_127 = {6{`RANDOM}};
  cache_data_124 = _RAND_127[184:0];
  _RAND_128 = {6{`RANDOM}};
  cache_data_125 = _RAND_128[184:0];
  _RAND_129 = {6{`RANDOM}};
  cache_data_126 = _RAND_129[184:0];
  _RAND_130 = {6{`RANDOM}};
  cache_data_127 = _RAND_130[184:0];
  _RAND_131 = {6{`RANDOM}};
  cache_data_128 = _RAND_131[184:0];
  _RAND_132 = {6{`RANDOM}};
  cache_data_129 = _RAND_132[184:0];
  _RAND_133 = {6{`RANDOM}};
  cache_data_130 = _RAND_133[184:0];
  _RAND_134 = {6{`RANDOM}};
  cache_data_131 = _RAND_134[184:0];
  _RAND_135 = {6{`RANDOM}};
  cache_data_132 = _RAND_135[184:0];
  _RAND_136 = {6{`RANDOM}};
  cache_data_133 = _RAND_136[184:0];
  _RAND_137 = {6{`RANDOM}};
  cache_data_134 = _RAND_137[184:0];
  _RAND_138 = {6{`RANDOM}};
  cache_data_135 = _RAND_138[184:0];
  _RAND_139 = {6{`RANDOM}};
  cache_data_136 = _RAND_139[184:0];
  _RAND_140 = {6{`RANDOM}};
  cache_data_137 = _RAND_140[184:0];
  _RAND_141 = {6{`RANDOM}};
  cache_data_138 = _RAND_141[184:0];
  _RAND_142 = {6{`RANDOM}};
  cache_data_139 = _RAND_142[184:0];
  _RAND_143 = {6{`RANDOM}};
  cache_data_140 = _RAND_143[184:0];
  _RAND_144 = {6{`RANDOM}};
  cache_data_141 = _RAND_144[184:0];
  _RAND_145 = {6{`RANDOM}};
  cache_data_142 = _RAND_145[184:0];
  _RAND_146 = {6{`RANDOM}};
  cache_data_143 = _RAND_146[184:0];
  _RAND_147 = {6{`RANDOM}};
  cache_data_144 = _RAND_147[184:0];
  _RAND_148 = {6{`RANDOM}};
  cache_data_145 = _RAND_148[184:0];
  _RAND_149 = {6{`RANDOM}};
  cache_data_146 = _RAND_149[184:0];
  _RAND_150 = {6{`RANDOM}};
  cache_data_147 = _RAND_150[184:0];
  _RAND_151 = {6{`RANDOM}};
  cache_data_148 = _RAND_151[184:0];
  _RAND_152 = {6{`RANDOM}};
  cache_data_149 = _RAND_152[184:0];
  _RAND_153 = {6{`RANDOM}};
  cache_data_150 = _RAND_153[184:0];
  _RAND_154 = {6{`RANDOM}};
  cache_data_151 = _RAND_154[184:0];
  _RAND_155 = {6{`RANDOM}};
  cache_data_152 = _RAND_155[184:0];
  _RAND_156 = {6{`RANDOM}};
  cache_data_153 = _RAND_156[184:0];
  _RAND_157 = {6{`RANDOM}};
  cache_data_154 = _RAND_157[184:0];
  _RAND_158 = {6{`RANDOM}};
  cache_data_155 = _RAND_158[184:0];
  _RAND_159 = {6{`RANDOM}};
  cache_data_156 = _RAND_159[184:0];
  _RAND_160 = {6{`RANDOM}};
  cache_data_157 = _RAND_160[184:0];
  _RAND_161 = {6{`RANDOM}};
  cache_data_158 = _RAND_161[184:0];
  _RAND_162 = {6{`RANDOM}};
  cache_data_159 = _RAND_162[184:0];
  _RAND_163 = {6{`RANDOM}};
  cache_data_160 = _RAND_163[184:0];
  _RAND_164 = {6{`RANDOM}};
  cache_data_161 = _RAND_164[184:0];
  _RAND_165 = {6{`RANDOM}};
  cache_data_162 = _RAND_165[184:0];
  _RAND_166 = {6{`RANDOM}};
  cache_data_163 = _RAND_166[184:0];
  _RAND_167 = {6{`RANDOM}};
  cache_data_164 = _RAND_167[184:0];
  _RAND_168 = {6{`RANDOM}};
  cache_data_165 = _RAND_168[184:0];
  _RAND_169 = {6{`RANDOM}};
  cache_data_166 = _RAND_169[184:0];
  _RAND_170 = {6{`RANDOM}};
  cache_data_167 = _RAND_170[184:0];
  _RAND_171 = {6{`RANDOM}};
  cache_data_168 = _RAND_171[184:0];
  _RAND_172 = {6{`RANDOM}};
  cache_data_169 = _RAND_172[184:0];
  _RAND_173 = {6{`RANDOM}};
  cache_data_170 = _RAND_173[184:0];
  _RAND_174 = {6{`RANDOM}};
  cache_data_171 = _RAND_174[184:0];
  _RAND_175 = {6{`RANDOM}};
  cache_data_172 = _RAND_175[184:0];
  _RAND_176 = {6{`RANDOM}};
  cache_data_173 = _RAND_176[184:0];
  _RAND_177 = {6{`RANDOM}};
  cache_data_174 = _RAND_177[184:0];
  _RAND_178 = {6{`RANDOM}};
  cache_data_175 = _RAND_178[184:0];
  _RAND_179 = {6{`RANDOM}};
  cache_data_176 = _RAND_179[184:0];
  _RAND_180 = {6{`RANDOM}};
  cache_data_177 = _RAND_180[184:0];
  _RAND_181 = {6{`RANDOM}};
  cache_data_178 = _RAND_181[184:0];
  _RAND_182 = {6{`RANDOM}};
  cache_data_179 = _RAND_182[184:0];
  _RAND_183 = {6{`RANDOM}};
  cache_data_180 = _RAND_183[184:0];
  _RAND_184 = {6{`RANDOM}};
  cache_data_181 = _RAND_184[184:0];
  _RAND_185 = {6{`RANDOM}};
  cache_data_182 = _RAND_185[184:0];
  _RAND_186 = {6{`RANDOM}};
  cache_data_183 = _RAND_186[184:0];
  _RAND_187 = {6{`RANDOM}};
  cache_data_184 = _RAND_187[184:0];
  _RAND_188 = {6{`RANDOM}};
  cache_data_185 = _RAND_188[184:0];
  _RAND_189 = {6{`RANDOM}};
  cache_data_186 = _RAND_189[184:0];
  _RAND_190 = {6{`RANDOM}};
  cache_data_187 = _RAND_190[184:0];
  _RAND_191 = {6{`RANDOM}};
  cache_data_188 = _RAND_191[184:0];
  _RAND_192 = {6{`RANDOM}};
  cache_data_189 = _RAND_192[184:0];
  _RAND_193 = {6{`RANDOM}};
  cache_data_190 = _RAND_193[184:0];
  _RAND_194 = {6{`RANDOM}};
  cache_data_191 = _RAND_194[184:0];
  _RAND_195 = {6{`RANDOM}};
  cache_data_192 = _RAND_195[184:0];
  _RAND_196 = {6{`RANDOM}};
  cache_data_193 = _RAND_196[184:0];
  _RAND_197 = {6{`RANDOM}};
  cache_data_194 = _RAND_197[184:0];
  _RAND_198 = {6{`RANDOM}};
  cache_data_195 = _RAND_198[184:0];
  _RAND_199 = {6{`RANDOM}};
  cache_data_196 = _RAND_199[184:0];
  _RAND_200 = {6{`RANDOM}};
  cache_data_197 = _RAND_200[184:0];
  _RAND_201 = {6{`RANDOM}};
  cache_data_198 = _RAND_201[184:0];
  _RAND_202 = {6{`RANDOM}};
  cache_data_199 = _RAND_202[184:0];
  _RAND_203 = {6{`RANDOM}};
  cache_data_200 = _RAND_203[184:0];
  _RAND_204 = {6{`RANDOM}};
  cache_data_201 = _RAND_204[184:0];
  _RAND_205 = {6{`RANDOM}};
  cache_data_202 = _RAND_205[184:0];
  _RAND_206 = {6{`RANDOM}};
  cache_data_203 = _RAND_206[184:0];
  _RAND_207 = {6{`RANDOM}};
  cache_data_204 = _RAND_207[184:0];
  _RAND_208 = {6{`RANDOM}};
  cache_data_205 = _RAND_208[184:0];
  _RAND_209 = {6{`RANDOM}};
  cache_data_206 = _RAND_209[184:0];
  _RAND_210 = {6{`RANDOM}};
  cache_data_207 = _RAND_210[184:0];
  _RAND_211 = {6{`RANDOM}};
  cache_data_208 = _RAND_211[184:0];
  _RAND_212 = {6{`RANDOM}};
  cache_data_209 = _RAND_212[184:0];
  _RAND_213 = {6{`RANDOM}};
  cache_data_210 = _RAND_213[184:0];
  _RAND_214 = {6{`RANDOM}};
  cache_data_211 = _RAND_214[184:0];
  _RAND_215 = {6{`RANDOM}};
  cache_data_212 = _RAND_215[184:0];
  _RAND_216 = {6{`RANDOM}};
  cache_data_213 = _RAND_216[184:0];
  _RAND_217 = {6{`RANDOM}};
  cache_data_214 = _RAND_217[184:0];
  _RAND_218 = {6{`RANDOM}};
  cache_data_215 = _RAND_218[184:0];
  _RAND_219 = {6{`RANDOM}};
  cache_data_216 = _RAND_219[184:0];
  _RAND_220 = {6{`RANDOM}};
  cache_data_217 = _RAND_220[184:0];
  _RAND_221 = {6{`RANDOM}};
  cache_data_218 = _RAND_221[184:0];
  _RAND_222 = {6{`RANDOM}};
  cache_data_219 = _RAND_222[184:0];
  _RAND_223 = {6{`RANDOM}};
  cache_data_220 = _RAND_223[184:0];
  _RAND_224 = {6{`RANDOM}};
  cache_data_221 = _RAND_224[184:0];
  _RAND_225 = {6{`RANDOM}};
  cache_data_222 = _RAND_225[184:0];
  _RAND_226 = {6{`RANDOM}};
  cache_data_223 = _RAND_226[184:0];
  _RAND_227 = {6{`RANDOM}};
  cache_data_224 = _RAND_227[184:0];
  _RAND_228 = {6{`RANDOM}};
  cache_data_225 = _RAND_228[184:0];
  _RAND_229 = {6{`RANDOM}};
  cache_data_226 = _RAND_229[184:0];
  _RAND_230 = {6{`RANDOM}};
  cache_data_227 = _RAND_230[184:0];
  _RAND_231 = {6{`RANDOM}};
  cache_data_228 = _RAND_231[184:0];
  _RAND_232 = {6{`RANDOM}};
  cache_data_229 = _RAND_232[184:0];
  _RAND_233 = {6{`RANDOM}};
  cache_data_230 = _RAND_233[184:0];
  _RAND_234 = {6{`RANDOM}};
  cache_data_231 = _RAND_234[184:0];
  _RAND_235 = {6{`RANDOM}};
  cache_data_232 = _RAND_235[184:0];
  _RAND_236 = {6{`RANDOM}};
  cache_data_233 = _RAND_236[184:0];
  _RAND_237 = {6{`RANDOM}};
  cache_data_234 = _RAND_237[184:0];
  _RAND_238 = {6{`RANDOM}};
  cache_data_235 = _RAND_238[184:0];
  _RAND_239 = {6{`RANDOM}};
  cache_data_236 = _RAND_239[184:0];
  _RAND_240 = {6{`RANDOM}};
  cache_data_237 = _RAND_240[184:0];
  _RAND_241 = {6{`RANDOM}};
  cache_data_238 = _RAND_241[184:0];
  _RAND_242 = {6{`RANDOM}};
  cache_data_239 = _RAND_242[184:0];
  _RAND_243 = {6{`RANDOM}};
  cache_data_240 = _RAND_243[184:0];
  _RAND_244 = {6{`RANDOM}};
  cache_data_241 = _RAND_244[184:0];
  _RAND_245 = {6{`RANDOM}};
  cache_data_242 = _RAND_245[184:0];
  _RAND_246 = {6{`RANDOM}};
  cache_data_243 = _RAND_246[184:0];
  _RAND_247 = {6{`RANDOM}};
  cache_data_244 = _RAND_247[184:0];
  _RAND_248 = {6{`RANDOM}};
  cache_data_245 = _RAND_248[184:0];
  _RAND_249 = {6{`RANDOM}};
  cache_data_246 = _RAND_249[184:0];
  _RAND_250 = {6{`RANDOM}};
  cache_data_247 = _RAND_250[184:0];
  _RAND_251 = {6{`RANDOM}};
  cache_data_248 = _RAND_251[184:0];
  _RAND_252 = {6{`RANDOM}};
  cache_data_249 = _RAND_252[184:0];
  _RAND_253 = {6{`RANDOM}};
  cache_data_250 = _RAND_253[184:0];
  _RAND_254 = {6{`RANDOM}};
  cache_data_251 = _RAND_254[184:0];
  _RAND_255 = {6{`RANDOM}};
  cache_data_252 = _RAND_255[184:0];
  _RAND_256 = {6{`RANDOM}};
  cache_data_253 = _RAND_256[184:0];
  _RAND_257 = {6{`RANDOM}};
  cache_data_254 = _RAND_257[184:0];
  _RAND_258 = {6{`RANDOM}};
  cache_data_255 = _RAND_258[184:0];
  _RAND_259 = {6{`RANDOM}};
  cache_data_256 = _RAND_259[184:0];
  _RAND_260 = {6{`RANDOM}};
  cache_data_257 = _RAND_260[184:0];
  _RAND_261 = {6{`RANDOM}};
  cache_data_258 = _RAND_261[184:0];
  _RAND_262 = {6{`RANDOM}};
  cache_data_259 = _RAND_262[184:0];
  _RAND_263 = {6{`RANDOM}};
  cache_data_260 = _RAND_263[184:0];
  _RAND_264 = {6{`RANDOM}};
  cache_data_261 = _RAND_264[184:0];
  _RAND_265 = {6{`RANDOM}};
  cache_data_262 = _RAND_265[184:0];
  _RAND_266 = {6{`RANDOM}};
  cache_data_263 = _RAND_266[184:0];
  _RAND_267 = {6{`RANDOM}};
  cache_data_264 = _RAND_267[184:0];
  _RAND_268 = {6{`RANDOM}};
  cache_data_265 = _RAND_268[184:0];
  _RAND_269 = {6{`RANDOM}};
  cache_data_266 = _RAND_269[184:0];
  _RAND_270 = {6{`RANDOM}};
  cache_data_267 = _RAND_270[184:0];
  _RAND_271 = {6{`RANDOM}};
  cache_data_268 = _RAND_271[184:0];
  _RAND_272 = {6{`RANDOM}};
  cache_data_269 = _RAND_272[184:0];
  _RAND_273 = {6{`RANDOM}};
  cache_data_270 = _RAND_273[184:0];
  _RAND_274 = {6{`RANDOM}};
  cache_data_271 = _RAND_274[184:0];
  _RAND_275 = {6{`RANDOM}};
  cache_data_272 = _RAND_275[184:0];
  _RAND_276 = {6{`RANDOM}};
  cache_data_273 = _RAND_276[184:0];
  _RAND_277 = {6{`RANDOM}};
  cache_data_274 = _RAND_277[184:0];
  _RAND_278 = {6{`RANDOM}};
  cache_data_275 = _RAND_278[184:0];
  _RAND_279 = {6{`RANDOM}};
  cache_data_276 = _RAND_279[184:0];
  _RAND_280 = {6{`RANDOM}};
  cache_data_277 = _RAND_280[184:0];
  _RAND_281 = {6{`RANDOM}};
  cache_data_278 = _RAND_281[184:0];
  _RAND_282 = {6{`RANDOM}};
  cache_data_279 = _RAND_282[184:0];
  _RAND_283 = {6{`RANDOM}};
  cache_data_280 = _RAND_283[184:0];
  _RAND_284 = {6{`RANDOM}};
  cache_data_281 = _RAND_284[184:0];
  _RAND_285 = {6{`RANDOM}};
  cache_data_282 = _RAND_285[184:0];
  _RAND_286 = {6{`RANDOM}};
  cache_data_283 = _RAND_286[184:0];
  _RAND_287 = {6{`RANDOM}};
  cache_data_284 = _RAND_287[184:0];
  _RAND_288 = {6{`RANDOM}};
  cache_data_285 = _RAND_288[184:0];
  _RAND_289 = {6{`RANDOM}};
  cache_data_286 = _RAND_289[184:0];
  _RAND_290 = {6{`RANDOM}};
  cache_data_287 = _RAND_290[184:0];
  _RAND_291 = {6{`RANDOM}};
  cache_data_288 = _RAND_291[184:0];
  _RAND_292 = {6{`RANDOM}};
  cache_data_289 = _RAND_292[184:0];
  _RAND_293 = {6{`RANDOM}};
  cache_data_290 = _RAND_293[184:0];
  _RAND_294 = {6{`RANDOM}};
  cache_data_291 = _RAND_294[184:0];
  _RAND_295 = {6{`RANDOM}};
  cache_data_292 = _RAND_295[184:0];
  _RAND_296 = {6{`RANDOM}};
  cache_data_293 = _RAND_296[184:0];
  _RAND_297 = {6{`RANDOM}};
  cache_data_294 = _RAND_297[184:0];
  _RAND_298 = {6{`RANDOM}};
  cache_data_295 = _RAND_298[184:0];
  _RAND_299 = {6{`RANDOM}};
  cache_data_296 = _RAND_299[184:0];
  _RAND_300 = {6{`RANDOM}};
  cache_data_297 = _RAND_300[184:0];
  _RAND_301 = {6{`RANDOM}};
  cache_data_298 = _RAND_301[184:0];
  _RAND_302 = {6{`RANDOM}};
  cache_data_299 = _RAND_302[184:0];
  _RAND_303 = {6{`RANDOM}};
  cache_data_300 = _RAND_303[184:0];
  _RAND_304 = {6{`RANDOM}};
  cache_data_301 = _RAND_304[184:0];
  _RAND_305 = {6{`RANDOM}};
  cache_data_302 = _RAND_305[184:0];
  _RAND_306 = {6{`RANDOM}};
  cache_data_303 = _RAND_306[184:0];
  _RAND_307 = {6{`RANDOM}};
  cache_data_304 = _RAND_307[184:0];
  _RAND_308 = {6{`RANDOM}};
  cache_data_305 = _RAND_308[184:0];
  _RAND_309 = {6{`RANDOM}};
  cache_data_306 = _RAND_309[184:0];
  _RAND_310 = {6{`RANDOM}};
  cache_data_307 = _RAND_310[184:0];
  _RAND_311 = {6{`RANDOM}};
  cache_data_308 = _RAND_311[184:0];
  _RAND_312 = {6{`RANDOM}};
  cache_data_309 = _RAND_312[184:0];
  _RAND_313 = {6{`RANDOM}};
  cache_data_310 = _RAND_313[184:0];
  _RAND_314 = {6{`RANDOM}};
  cache_data_311 = _RAND_314[184:0];
  _RAND_315 = {6{`RANDOM}};
  cache_data_312 = _RAND_315[184:0];
  _RAND_316 = {6{`RANDOM}};
  cache_data_313 = _RAND_316[184:0];
  _RAND_317 = {6{`RANDOM}};
  cache_data_314 = _RAND_317[184:0];
  _RAND_318 = {6{`RANDOM}};
  cache_data_315 = _RAND_318[184:0];
  _RAND_319 = {6{`RANDOM}};
  cache_data_316 = _RAND_319[184:0];
  _RAND_320 = {6{`RANDOM}};
  cache_data_317 = _RAND_320[184:0];
  _RAND_321 = {6{`RANDOM}};
  cache_data_318 = _RAND_321[184:0];
  _RAND_322 = {6{`RANDOM}};
  cache_data_319 = _RAND_322[184:0];
  _RAND_323 = {6{`RANDOM}};
  cache_data_320 = _RAND_323[184:0];
  _RAND_324 = {6{`RANDOM}};
  cache_data_321 = _RAND_324[184:0];
  _RAND_325 = {6{`RANDOM}};
  cache_data_322 = _RAND_325[184:0];
  _RAND_326 = {6{`RANDOM}};
  cache_data_323 = _RAND_326[184:0];
  _RAND_327 = {6{`RANDOM}};
  cache_data_324 = _RAND_327[184:0];
  _RAND_328 = {6{`RANDOM}};
  cache_data_325 = _RAND_328[184:0];
  _RAND_329 = {6{`RANDOM}};
  cache_data_326 = _RAND_329[184:0];
  _RAND_330 = {6{`RANDOM}};
  cache_data_327 = _RAND_330[184:0];
  _RAND_331 = {6{`RANDOM}};
  cache_data_328 = _RAND_331[184:0];
  _RAND_332 = {6{`RANDOM}};
  cache_data_329 = _RAND_332[184:0];
  _RAND_333 = {6{`RANDOM}};
  cache_data_330 = _RAND_333[184:0];
  _RAND_334 = {6{`RANDOM}};
  cache_data_331 = _RAND_334[184:0];
  _RAND_335 = {6{`RANDOM}};
  cache_data_332 = _RAND_335[184:0];
  _RAND_336 = {6{`RANDOM}};
  cache_data_333 = _RAND_336[184:0];
  _RAND_337 = {6{`RANDOM}};
  cache_data_334 = _RAND_337[184:0];
  _RAND_338 = {6{`RANDOM}};
  cache_data_335 = _RAND_338[184:0];
  _RAND_339 = {6{`RANDOM}};
  cache_data_336 = _RAND_339[184:0];
  _RAND_340 = {6{`RANDOM}};
  cache_data_337 = _RAND_340[184:0];
  _RAND_341 = {6{`RANDOM}};
  cache_data_338 = _RAND_341[184:0];
  _RAND_342 = {6{`RANDOM}};
  cache_data_339 = _RAND_342[184:0];
  _RAND_343 = {6{`RANDOM}};
  cache_data_340 = _RAND_343[184:0];
  _RAND_344 = {6{`RANDOM}};
  cache_data_341 = _RAND_344[184:0];
  _RAND_345 = {6{`RANDOM}};
  cache_data_342 = _RAND_345[184:0];
  _RAND_346 = {6{`RANDOM}};
  cache_data_343 = _RAND_346[184:0];
  _RAND_347 = {6{`RANDOM}};
  cache_data_344 = _RAND_347[184:0];
  _RAND_348 = {6{`RANDOM}};
  cache_data_345 = _RAND_348[184:0];
  _RAND_349 = {6{`RANDOM}};
  cache_data_346 = _RAND_349[184:0];
  _RAND_350 = {6{`RANDOM}};
  cache_data_347 = _RAND_350[184:0];
  _RAND_351 = {6{`RANDOM}};
  cache_data_348 = _RAND_351[184:0];
  _RAND_352 = {6{`RANDOM}};
  cache_data_349 = _RAND_352[184:0];
  _RAND_353 = {6{`RANDOM}};
  cache_data_350 = _RAND_353[184:0];
  _RAND_354 = {6{`RANDOM}};
  cache_data_351 = _RAND_354[184:0];
  _RAND_355 = {6{`RANDOM}};
  cache_data_352 = _RAND_355[184:0];
  _RAND_356 = {6{`RANDOM}};
  cache_data_353 = _RAND_356[184:0];
  _RAND_357 = {6{`RANDOM}};
  cache_data_354 = _RAND_357[184:0];
  _RAND_358 = {6{`RANDOM}};
  cache_data_355 = _RAND_358[184:0];
  _RAND_359 = {6{`RANDOM}};
  cache_data_356 = _RAND_359[184:0];
  _RAND_360 = {6{`RANDOM}};
  cache_data_357 = _RAND_360[184:0];
  _RAND_361 = {6{`RANDOM}};
  cache_data_358 = _RAND_361[184:0];
  _RAND_362 = {6{`RANDOM}};
  cache_data_359 = _RAND_362[184:0];
  _RAND_363 = {6{`RANDOM}};
  cache_data_360 = _RAND_363[184:0];
  _RAND_364 = {6{`RANDOM}};
  cache_data_361 = _RAND_364[184:0];
  _RAND_365 = {6{`RANDOM}};
  cache_data_362 = _RAND_365[184:0];
  _RAND_366 = {6{`RANDOM}};
  cache_data_363 = _RAND_366[184:0];
  _RAND_367 = {6{`RANDOM}};
  cache_data_364 = _RAND_367[184:0];
  _RAND_368 = {6{`RANDOM}};
  cache_data_365 = _RAND_368[184:0];
  _RAND_369 = {6{`RANDOM}};
  cache_data_366 = _RAND_369[184:0];
  _RAND_370 = {6{`RANDOM}};
  cache_data_367 = _RAND_370[184:0];
  _RAND_371 = {6{`RANDOM}};
  cache_data_368 = _RAND_371[184:0];
  _RAND_372 = {6{`RANDOM}};
  cache_data_369 = _RAND_372[184:0];
  _RAND_373 = {6{`RANDOM}};
  cache_data_370 = _RAND_373[184:0];
  _RAND_374 = {6{`RANDOM}};
  cache_data_371 = _RAND_374[184:0];
  _RAND_375 = {6{`RANDOM}};
  cache_data_372 = _RAND_375[184:0];
  _RAND_376 = {6{`RANDOM}};
  cache_data_373 = _RAND_376[184:0];
  _RAND_377 = {6{`RANDOM}};
  cache_data_374 = _RAND_377[184:0];
  _RAND_378 = {6{`RANDOM}};
  cache_data_375 = _RAND_378[184:0];
  _RAND_379 = {6{`RANDOM}};
  cache_data_376 = _RAND_379[184:0];
  _RAND_380 = {6{`RANDOM}};
  cache_data_377 = _RAND_380[184:0];
  _RAND_381 = {6{`RANDOM}};
  cache_data_378 = _RAND_381[184:0];
  _RAND_382 = {6{`RANDOM}};
  cache_data_379 = _RAND_382[184:0];
  _RAND_383 = {6{`RANDOM}};
  cache_data_380 = _RAND_383[184:0];
  _RAND_384 = {6{`RANDOM}};
  cache_data_381 = _RAND_384[184:0];
  _RAND_385 = {6{`RANDOM}};
  cache_data_382 = _RAND_385[184:0];
  _RAND_386 = {6{`RANDOM}};
  cache_data_383 = _RAND_386[184:0];
  _RAND_387 = {6{`RANDOM}};
  cache_data_384 = _RAND_387[184:0];
  _RAND_388 = {6{`RANDOM}};
  cache_data_385 = _RAND_388[184:0];
  _RAND_389 = {6{`RANDOM}};
  cache_data_386 = _RAND_389[184:0];
  _RAND_390 = {6{`RANDOM}};
  cache_data_387 = _RAND_390[184:0];
  _RAND_391 = {6{`RANDOM}};
  cache_data_388 = _RAND_391[184:0];
  _RAND_392 = {6{`RANDOM}};
  cache_data_389 = _RAND_392[184:0];
  _RAND_393 = {6{`RANDOM}};
  cache_data_390 = _RAND_393[184:0];
  _RAND_394 = {6{`RANDOM}};
  cache_data_391 = _RAND_394[184:0];
  _RAND_395 = {6{`RANDOM}};
  cache_data_392 = _RAND_395[184:0];
  _RAND_396 = {6{`RANDOM}};
  cache_data_393 = _RAND_396[184:0];
  _RAND_397 = {6{`RANDOM}};
  cache_data_394 = _RAND_397[184:0];
  _RAND_398 = {6{`RANDOM}};
  cache_data_395 = _RAND_398[184:0];
  _RAND_399 = {6{`RANDOM}};
  cache_data_396 = _RAND_399[184:0];
  _RAND_400 = {6{`RANDOM}};
  cache_data_397 = _RAND_400[184:0];
  _RAND_401 = {6{`RANDOM}};
  cache_data_398 = _RAND_401[184:0];
  _RAND_402 = {6{`RANDOM}};
  cache_data_399 = _RAND_402[184:0];
  _RAND_403 = {6{`RANDOM}};
  cache_data_400 = _RAND_403[184:0];
  _RAND_404 = {6{`RANDOM}};
  cache_data_401 = _RAND_404[184:0];
  _RAND_405 = {6{`RANDOM}};
  cache_data_402 = _RAND_405[184:0];
  _RAND_406 = {6{`RANDOM}};
  cache_data_403 = _RAND_406[184:0];
  _RAND_407 = {6{`RANDOM}};
  cache_data_404 = _RAND_407[184:0];
  _RAND_408 = {6{`RANDOM}};
  cache_data_405 = _RAND_408[184:0];
  _RAND_409 = {6{`RANDOM}};
  cache_data_406 = _RAND_409[184:0];
  _RAND_410 = {6{`RANDOM}};
  cache_data_407 = _RAND_410[184:0];
  _RAND_411 = {6{`RANDOM}};
  cache_data_408 = _RAND_411[184:0];
  _RAND_412 = {6{`RANDOM}};
  cache_data_409 = _RAND_412[184:0];
  _RAND_413 = {6{`RANDOM}};
  cache_data_410 = _RAND_413[184:0];
  _RAND_414 = {6{`RANDOM}};
  cache_data_411 = _RAND_414[184:0];
  _RAND_415 = {6{`RANDOM}};
  cache_data_412 = _RAND_415[184:0];
  _RAND_416 = {6{`RANDOM}};
  cache_data_413 = _RAND_416[184:0];
  _RAND_417 = {6{`RANDOM}};
  cache_data_414 = _RAND_417[184:0];
  _RAND_418 = {6{`RANDOM}};
  cache_data_415 = _RAND_418[184:0];
  _RAND_419 = {6{`RANDOM}};
  cache_data_416 = _RAND_419[184:0];
  _RAND_420 = {6{`RANDOM}};
  cache_data_417 = _RAND_420[184:0];
  _RAND_421 = {6{`RANDOM}};
  cache_data_418 = _RAND_421[184:0];
  _RAND_422 = {6{`RANDOM}};
  cache_data_419 = _RAND_422[184:0];
  _RAND_423 = {6{`RANDOM}};
  cache_data_420 = _RAND_423[184:0];
  _RAND_424 = {6{`RANDOM}};
  cache_data_421 = _RAND_424[184:0];
  _RAND_425 = {6{`RANDOM}};
  cache_data_422 = _RAND_425[184:0];
  _RAND_426 = {6{`RANDOM}};
  cache_data_423 = _RAND_426[184:0];
  _RAND_427 = {6{`RANDOM}};
  cache_data_424 = _RAND_427[184:0];
  _RAND_428 = {6{`RANDOM}};
  cache_data_425 = _RAND_428[184:0];
  _RAND_429 = {6{`RANDOM}};
  cache_data_426 = _RAND_429[184:0];
  _RAND_430 = {6{`RANDOM}};
  cache_data_427 = _RAND_430[184:0];
  _RAND_431 = {6{`RANDOM}};
  cache_data_428 = _RAND_431[184:0];
  _RAND_432 = {6{`RANDOM}};
  cache_data_429 = _RAND_432[184:0];
  _RAND_433 = {6{`RANDOM}};
  cache_data_430 = _RAND_433[184:0];
  _RAND_434 = {6{`RANDOM}};
  cache_data_431 = _RAND_434[184:0];
  _RAND_435 = {6{`RANDOM}};
  cache_data_432 = _RAND_435[184:0];
  _RAND_436 = {6{`RANDOM}};
  cache_data_433 = _RAND_436[184:0];
  _RAND_437 = {6{`RANDOM}};
  cache_data_434 = _RAND_437[184:0];
  _RAND_438 = {6{`RANDOM}};
  cache_data_435 = _RAND_438[184:0];
  _RAND_439 = {6{`RANDOM}};
  cache_data_436 = _RAND_439[184:0];
  _RAND_440 = {6{`RANDOM}};
  cache_data_437 = _RAND_440[184:0];
  _RAND_441 = {6{`RANDOM}};
  cache_data_438 = _RAND_441[184:0];
  _RAND_442 = {6{`RANDOM}};
  cache_data_439 = _RAND_442[184:0];
  _RAND_443 = {6{`RANDOM}};
  cache_data_440 = _RAND_443[184:0];
  _RAND_444 = {6{`RANDOM}};
  cache_data_441 = _RAND_444[184:0];
  _RAND_445 = {6{`RANDOM}};
  cache_data_442 = _RAND_445[184:0];
  _RAND_446 = {6{`RANDOM}};
  cache_data_443 = _RAND_446[184:0];
  _RAND_447 = {6{`RANDOM}};
  cache_data_444 = _RAND_447[184:0];
  _RAND_448 = {6{`RANDOM}};
  cache_data_445 = _RAND_448[184:0];
  _RAND_449 = {6{`RANDOM}};
  cache_data_446 = _RAND_449[184:0];
  _RAND_450 = {6{`RANDOM}};
  cache_data_447 = _RAND_450[184:0];
  _RAND_451 = {6{`RANDOM}};
  cache_data_448 = _RAND_451[184:0];
  _RAND_452 = {6{`RANDOM}};
  cache_data_449 = _RAND_452[184:0];
  _RAND_453 = {6{`RANDOM}};
  cache_data_450 = _RAND_453[184:0];
  _RAND_454 = {6{`RANDOM}};
  cache_data_451 = _RAND_454[184:0];
  _RAND_455 = {6{`RANDOM}};
  cache_data_452 = _RAND_455[184:0];
  _RAND_456 = {6{`RANDOM}};
  cache_data_453 = _RAND_456[184:0];
  _RAND_457 = {6{`RANDOM}};
  cache_data_454 = _RAND_457[184:0];
  _RAND_458 = {6{`RANDOM}};
  cache_data_455 = _RAND_458[184:0];
  _RAND_459 = {6{`RANDOM}};
  cache_data_456 = _RAND_459[184:0];
  _RAND_460 = {6{`RANDOM}};
  cache_data_457 = _RAND_460[184:0];
  _RAND_461 = {6{`RANDOM}};
  cache_data_458 = _RAND_461[184:0];
  _RAND_462 = {6{`RANDOM}};
  cache_data_459 = _RAND_462[184:0];
  _RAND_463 = {6{`RANDOM}};
  cache_data_460 = _RAND_463[184:0];
  _RAND_464 = {6{`RANDOM}};
  cache_data_461 = _RAND_464[184:0];
  _RAND_465 = {6{`RANDOM}};
  cache_data_462 = _RAND_465[184:0];
  _RAND_466 = {6{`RANDOM}};
  cache_data_463 = _RAND_466[184:0];
  _RAND_467 = {6{`RANDOM}};
  cache_data_464 = _RAND_467[184:0];
  _RAND_468 = {6{`RANDOM}};
  cache_data_465 = _RAND_468[184:0];
  _RAND_469 = {6{`RANDOM}};
  cache_data_466 = _RAND_469[184:0];
  _RAND_470 = {6{`RANDOM}};
  cache_data_467 = _RAND_470[184:0];
  _RAND_471 = {6{`RANDOM}};
  cache_data_468 = _RAND_471[184:0];
  _RAND_472 = {6{`RANDOM}};
  cache_data_469 = _RAND_472[184:0];
  _RAND_473 = {6{`RANDOM}};
  cache_data_470 = _RAND_473[184:0];
  _RAND_474 = {6{`RANDOM}};
  cache_data_471 = _RAND_474[184:0];
  _RAND_475 = {6{`RANDOM}};
  cache_data_472 = _RAND_475[184:0];
  _RAND_476 = {6{`RANDOM}};
  cache_data_473 = _RAND_476[184:0];
  _RAND_477 = {6{`RANDOM}};
  cache_data_474 = _RAND_477[184:0];
  _RAND_478 = {6{`RANDOM}};
  cache_data_475 = _RAND_478[184:0];
  _RAND_479 = {6{`RANDOM}};
  cache_data_476 = _RAND_479[184:0];
  _RAND_480 = {6{`RANDOM}};
  cache_data_477 = _RAND_480[184:0];
  _RAND_481 = {6{`RANDOM}};
  cache_data_478 = _RAND_481[184:0];
  _RAND_482 = {6{`RANDOM}};
  cache_data_479 = _RAND_482[184:0];
  _RAND_483 = {6{`RANDOM}};
  cache_data_480 = _RAND_483[184:0];
  _RAND_484 = {6{`RANDOM}};
  cache_data_481 = _RAND_484[184:0];
  _RAND_485 = {6{`RANDOM}};
  cache_data_482 = _RAND_485[184:0];
  _RAND_486 = {6{`RANDOM}};
  cache_data_483 = _RAND_486[184:0];
  _RAND_487 = {6{`RANDOM}};
  cache_data_484 = _RAND_487[184:0];
  _RAND_488 = {6{`RANDOM}};
  cache_data_485 = _RAND_488[184:0];
  _RAND_489 = {6{`RANDOM}};
  cache_data_486 = _RAND_489[184:0];
  _RAND_490 = {6{`RANDOM}};
  cache_data_487 = _RAND_490[184:0];
  _RAND_491 = {6{`RANDOM}};
  cache_data_488 = _RAND_491[184:0];
  _RAND_492 = {6{`RANDOM}};
  cache_data_489 = _RAND_492[184:0];
  _RAND_493 = {6{`RANDOM}};
  cache_data_490 = _RAND_493[184:0];
  _RAND_494 = {6{`RANDOM}};
  cache_data_491 = _RAND_494[184:0];
  _RAND_495 = {6{`RANDOM}};
  cache_data_492 = _RAND_495[184:0];
  _RAND_496 = {6{`RANDOM}};
  cache_data_493 = _RAND_496[184:0];
  _RAND_497 = {6{`RANDOM}};
  cache_data_494 = _RAND_497[184:0];
  _RAND_498 = {6{`RANDOM}};
  cache_data_495 = _RAND_498[184:0];
  _RAND_499 = {6{`RANDOM}};
  cache_data_496 = _RAND_499[184:0];
  _RAND_500 = {6{`RANDOM}};
  cache_data_497 = _RAND_500[184:0];
  _RAND_501 = {6{`RANDOM}};
  cache_data_498 = _RAND_501[184:0];
  _RAND_502 = {6{`RANDOM}};
  cache_data_499 = _RAND_502[184:0];
  _RAND_503 = {6{`RANDOM}};
  cache_data_500 = _RAND_503[184:0];
  _RAND_504 = {6{`RANDOM}};
  cache_data_501 = _RAND_504[184:0];
  _RAND_505 = {6{`RANDOM}};
  cache_data_502 = _RAND_505[184:0];
  _RAND_506 = {6{`RANDOM}};
  cache_data_503 = _RAND_506[184:0];
  _RAND_507 = {6{`RANDOM}};
  cache_data_504 = _RAND_507[184:0];
  _RAND_508 = {6{`RANDOM}};
  cache_data_505 = _RAND_508[184:0];
  _RAND_509 = {6{`RANDOM}};
  cache_data_506 = _RAND_509[184:0];
  _RAND_510 = {6{`RANDOM}};
  cache_data_507 = _RAND_510[184:0];
  _RAND_511 = {6{`RANDOM}};
  cache_data_508 = _RAND_511[184:0];
  _RAND_512 = {6{`RANDOM}};
  cache_data_509 = _RAND_512[184:0];
  _RAND_513 = {6{`RANDOM}};
  cache_data_510 = _RAND_513[184:0];
  _RAND_514 = {6{`RANDOM}};
  cache_data_511 = _RAND_514[184:0];
  _RAND_515 = {6{`RANDOM}};
  cache_data_512 = _RAND_515[184:0];
  _RAND_516 = {6{`RANDOM}};
  cache_data_513 = _RAND_516[184:0];
  _RAND_517 = {6{`RANDOM}};
  cache_data_514 = _RAND_517[184:0];
  _RAND_518 = {6{`RANDOM}};
  cache_data_515 = _RAND_518[184:0];
  _RAND_519 = {6{`RANDOM}};
  cache_data_516 = _RAND_519[184:0];
  _RAND_520 = {6{`RANDOM}};
  cache_data_517 = _RAND_520[184:0];
  _RAND_521 = {6{`RANDOM}};
  cache_data_518 = _RAND_521[184:0];
  _RAND_522 = {6{`RANDOM}};
  cache_data_519 = _RAND_522[184:0];
  _RAND_523 = {6{`RANDOM}};
  cache_data_520 = _RAND_523[184:0];
  _RAND_524 = {6{`RANDOM}};
  cache_data_521 = _RAND_524[184:0];
  _RAND_525 = {6{`RANDOM}};
  cache_data_522 = _RAND_525[184:0];
  _RAND_526 = {6{`RANDOM}};
  cache_data_523 = _RAND_526[184:0];
  _RAND_527 = {6{`RANDOM}};
  cache_data_524 = _RAND_527[184:0];
  _RAND_528 = {6{`RANDOM}};
  cache_data_525 = _RAND_528[184:0];
  _RAND_529 = {6{`RANDOM}};
  cache_data_526 = _RAND_529[184:0];
  _RAND_530 = {6{`RANDOM}};
  cache_data_527 = _RAND_530[184:0];
  _RAND_531 = {6{`RANDOM}};
  cache_data_528 = _RAND_531[184:0];
  _RAND_532 = {6{`RANDOM}};
  cache_data_529 = _RAND_532[184:0];
  _RAND_533 = {6{`RANDOM}};
  cache_data_530 = _RAND_533[184:0];
  _RAND_534 = {6{`RANDOM}};
  cache_data_531 = _RAND_534[184:0];
  _RAND_535 = {6{`RANDOM}};
  cache_data_532 = _RAND_535[184:0];
  _RAND_536 = {6{`RANDOM}};
  cache_data_533 = _RAND_536[184:0];
  _RAND_537 = {6{`RANDOM}};
  cache_data_534 = _RAND_537[184:0];
  _RAND_538 = {6{`RANDOM}};
  cache_data_535 = _RAND_538[184:0];
  _RAND_539 = {6{`RANDOM}};
  cache_data_536 = _RAND_539[184:0];
  _RAND_540 = {6{`RANDOM}};
  cache_data_537 = _RAND_540[184:0];
  _RAND_541 = {6{`RANDOM}};
  cache_data_538 = _RAND_541[184:0];
  _RAND_542 = {6{`RANDOM}};
  cache_data_539 = _RAND_542[184:0];
  _RAND_543 = {6{`RANDOM}};
  cache_data_540 = _RAND_543[184:0];
  _RAND_544 = {6{`RANDOM}};
  cache_data_541 = _RAND_544[184:0];
  _RAND_545 = {6{`RANDOM}};
  cache_data_542 = _RAND_545[184:0];
  _RAND_546 = {6{`RANDOM}};
  cache_data_543 = _RAND_546[184:0];
  _RAND_547 = {6{`RANDOM}};
  cache_data_544 = _RAND_547[184:0];
  _RAND_548 = {6{`RANDOM}};
  cache_data_545 = _RAND_548[184:0];
  _RAND_549 = {6{`RANDOM}};
  cache_data_546 = _RAND_549[184:0];
  _RAND_550 = {6{`RANDOM}};
  cache_data_547 = _RAND_550[184:0];
  _RAND_551 = {6{`RANDOM}};
  cache_data_548 = _RAND_551[184:0];
  _RAND_552 = {6{`RANDOM}};
  cache_data_549 = _RAND_552[184:0];
  _RAND_553 = {6{`RANDOM}};
  cache_data_550 = _RAND_553[184:0];
  _RAND_554 = {6{`RANDOM}};
  cache_data_551 = _RAND_554[184:0];
  _RAND_555 = {6{`RANDOM}};
  cache_data_552 = _RAND_555[184:0];
  _RAND_556 = {6{`RANDOM}};
  cache_data_553 = _RAND_556[184:0];
  _RAND_557 = {6{`RANDOM}};
  cache_data_554 = _RAND_557[184:0];
  _RAND_558 = {6{`RANDOM}};
  cache_data_555 = _RAND_558[184:0];
  _RAND_559 = {6{`RANDOM}};
  cache_data_556 = _RAND_559[184:0];
  _RAND_560 = {6{`RANDOM}};
  cache_data_557 = _RAND_560[184:0];
  _RAND_561 = {6{`RANDOM}};
  cache_data_558 = _RAND_561[184:0];
  _RAND_562 = {6{`RANDOM}};
  cache_data_559 = _RAND_562[184:0];
  _RAND_563 = {6{`RANDOM}};
  cache_data_560 = _RAND_563[184:0];
  _RAND_564 = {6{`RANDOM}};
  cache_data_561 = _RAND_564[184:0];
  _RAND_565 = {6{`RANDOM}};
  cache_data_562 = _RAND_565[184:0];
  _RAND_566 = {6{`RANDOM}};
  cache_data_563 = _RAND_566[184:0];
  _RAND_567 = {6{`RANDOM}};
  cache_data_564 = _RAND_567[184:0];
  _RAND_568 = {6{`RANDOM}};
  cache_data_565 = _RAND_568[184:0];
  _RAND_569 = {6{`RANDOM}};
  cache_data_566 = _RAND_569[184:0];
  _RAND_570 = {6{`RANDOM}};
  cache_data_567 = _RAND_570[184:0];
  _RAND_571 = {6{`RANDOM}};
  cache_data_568 = _RAND_571[184:0];
  _RAND_572 = {6{`RANDOM}};
  cache_data_569 = _RAND_572[184:0];
  _RAND_573 = {6{`RANDOM}};
  cache_data_570 = _RAND_573[184:0];
  _RAND_574 = {6{`RANDOM}};
  cache_data_571 = _RAND_574[184:0];
  _RAND_575 = {6{`RANDOM}};
  cache_data_572 = _RAND_575[184:0];
  _RAND_576 = {6{`RANDOM}};
  cache_data_573 = _RAND_576[184:0];
  _RAND_577 = {6{`RANDOM}};
  cache_data_574 = _RAND_577[184:0];
  _RAND_578 = {6{`RANDOM}};
  cache_data_575 = _RAND_578[184:0];
  _RAND_579 = {6{`RANDOM}};
  cache_data_576 = _RAND_579[184:0];
  _RAND_580 = {6{`RANDOM}};
  cache_data_577 = _RAND_580[184:0];
  _RAND_581 = {6{`RANDOM}};
  cache_data_578 = _RAND_581[184:0];
  _RAND_582 = {6{`RANDOM}};
  cache_data_579 = _RAND_582[184:0];
  _RAND_583 = {6{`RANDOM}};
  cache_data_580 = _RAND_583[184:0];
  _RAND_584 = {6{`RANDOM}};
  cache_data_581 = _RAND_584[184:0];
  _RAND_585 = {6{`RANDOM}};
  cache_data_582 = _RAND_585[184:0];
  _RAND_586 = {6{`RANDOM}};
  cache_data_583 = _RAND_586[184:0];
  _RAND_587 = {6{`RANDOM}};
  cache_data_584 = _RAND_587[184:0];
  _RAND_588 = {6{`RANDOM}};
  cache_data_585 = _RAND_588[184:0];
  _RAND_589 = {6{`RANDOM}};
  cache_data_586 = _RAND_589[184:0];
  _RAND_590 = {6{`RANDOM}};
  cache_data_587 = _RAND_590[184:0];
  _RAND_591 = {6{`RANDOM}};
  cache_data_588 = _RAND_591[184:0];
  _RAND_592 = {6{`RANDOM}};
  cache_data_589 = _RAND_592[184:0];
  _RAND_593 = {6{`RANDOM}};
  cache_data_590 = _RAND_593[184:0];
  _RAND_594 = {6{`RANDOM}};
  cache_data_591 = _RAND_594[184:0];
  _RAND_595 = {6{`RANDOM}};
  cache_data_592 = _RAND_595[184:0];
  _RAND_596 = {6{`RANDOM}};
  cache_data_593 = _RAND_596[184:0];
  _RAND_597 = {6{`RANDOM}};
  cache_data_594 = _RAND_597[184:0];
  _RAND_598 = {6{`RANDOM}};
  cache_data_595 = _RAND_598[184:0];
  _RAND_599 = {6{`RANDOM}};
  cache_data_596 = _RAND_599[184:0];
  _RAND_600 = {6{`RANDOM}};
  cache_data_597 = _RAND_600[184:0];
  _RAND_601 = {6{`RANDOM}};
  cache_data_598 = _RAND_601[184:0];
  _RAND_602 = {6{`RANDOM}};
  cache_data_599 = _RAND_602[184:0];
  _RAND_603 = {6{`RANDOM}};
  cache_data_600 = _RAND_603[184:0];
  _RAND_604 = {6{`RANDOM}};
  cache_data_601 = _RAND_604[184:0];
  _RAND_605 = {6{`RANDOM}};
  cache_data_602 = _RAND_605[184:0];
  _RAND_606 = {6{`RANDOM}};
  cache_data_603 = _RAND_606[184:0];
  _RAND_607 = {6{`RANDOM}};
  cache_data_604 = _RAND_607[184:0];
  _RAND_608 = {6{`RANDOM}};
  cache_data_605 = _RAND_608[184:0];
  _RAND_609 = {6{`RANDOM}};
  cache_data_606 = _RAND_609[184:0];
  _RAND_610 = {6{`RANDOM}};
  cache_data_607 = _RAND_610[184:0];
  _RAND_611 = {6{`RANDOM}};
  cache_data_608 = _RAND_611[184:0];
  _RAND_612 = {6{`RANDOM}};
  cache_data_609 = _RAND_612[184:0];
  _RAND_613 = {6{`RANDOM}};
  cache_data_610 = _RAND_613[184:0];
  _RAND_614 = {6{`RANDOM}};
  cache_data_611 = _RAND_614[184:0];
  _RAND_615 = {6{`RANDOM}};
  cache_data_612 = _RAND_615[184:0];
  _RAND_616 = {6{`RANDOM}};
  cache_data_613 = _RAND_616[184:0];
  _RAND_617 = {6{`RANDOM}};
  cache_data_614 = _RAND_617[184:0];
  _RAND_618 = {6{`RANDOM}};
  cache_data_615 = _RAND_618[184:0];
  _RAND_619 = {6{`RANDOM}};
  cache_data_616 = _RAND_619[184:0];
  _RAND_620 = {6{`RANDOM}};
  cache_data_617 = _RAND_620[184:0];
  _RAND_621 = {6{`RANDOM}};
  cache_data_618 = _RAND_621[184:0];
  _RAND_622 = {6{`RANDOM}};
  cache_data_619 = _RAND_622[184:0];
  _RAND_623 = {6{`RANDOM}};
  cache_data_620 = _RAND_623[184:0];
  _RAND_624 = {6{`RANDOM}};
  cache_data_621 = _RAND_624[184:0];
  _RAND_625 = {6{`RANDOM}};
  cache_data_622 = _RAND_625[184:0];
  _RAND_626 = {6{`RANDOM}};
  cache_data_623 = _RAND_626[184:0];
  _RAND_627 = {6{`RANDOM}};
  cache_data_624 = _RAND_627[184:0];
  _RAND_628 = {6{`RANDOM}};
  cache_data_625 = _RAND_628[184:0];
  _RAND_629 = {6{`RANDOM}};
  cache_data_626 = _RAND_629[184:0];
  _RAND_630 = {6{`RANDOM}};
  cache_data_627 = _RAND_630[184:0];
  _RAND_631 = {6{`RANDOM}};
  cache_data_628 = _RAND_631[184:0];
  _RAND_632 = {6{`RANDOM}};
  cache_data_629 = _RAND_632[184:0];
  _RAND_633 = {6{`RANDOM}};
  cache_data_630 = _RAND_633[184:0];
  _RAND_634 = {6{`RANDOM}};
  cache_data_631 = _RAND_634[184:0];
  _RAND_635 = {6{`RANDOM}};
  cache_data_632 = _RAND_635[184:0];
  _RAND_636 = {6{`RANDOM}};
  cache_data_633 = _RAND_636[184:0];
  _RAND_637 = {6{`RANDOM}};
  cache_data_634 = _RAND_637[184:0];
  _RAND_638 = {6{`RANDOM}};
  cache_data_635 = _RAND_638[184:0];
  _RAND_639 = {6{`RANDOM}};
  cache_data_636 = _RAND_639[184:0];
  _RAND_640 = {6{`RANDOM}};
  cache_data_637 = _RAND_640[184:0];
  _RAND_641 = {6{`RANDOM}};
  cache_data_638 = _RAND_641[184:0];
  _RAND_642 = {6{`RANDOM}};
  cache_data_639 = _RAND_642[184:0];
  _RAND_643 = {6{`RANDOM}};
  cache_data_640 = _RAND_643[184:0];
  _RAND_644 = {6{`RANDOM}};
  cache_data_641 = _RAND_644[184:0];
  _RAND_645 = {6{`RANDOM}};
  cache_data_642 = _RAND_645[184:0];
  _RAND_646 = {6{`RANDOM}};
  cache_data_643 = _RAND_646[184:0];
  _RAND_647 = {6{`RANDOM}};
  cache_data_644 = _RAND_647[184:0];
  _RAND_648 = {6{`RANDOM}};
  cache_data_645 = _RAND_648[184:0];
  _RAND_649 = {6{`RANDOM}};
  cache_data_646 = _RAND_649[184:0];
  _RAND_650 = {6{`RANDOM}};
  cache_data_647 = _RAND_650[184:0];
  _RAND_651 = {6{`RANDOM}};
  cache_data_648 = _RAND_651[184:0];
  _RAND_652 = {6{`RANDOM}};
  cache_data_649 = _RAND_652[184:0];
  _RAND_653 = {6{`RANDOM}};
  cache_data_650 = _RAND_653[184:0];
  _RAND_654 = {6{`RANDOM}};
  cache_data_651 = _RAND_654[184:0];
  _RAND_655 = {6{`RANDOM}};
  cache_data_652 = _RAND_655[184:0];
  _RAND_656 = {6{`RANDOM}};
  cache_data_653 = _RAND_656[184:0];
  _RAND_657 = {6{`RANDOM}};
  cache_data_654 = _RAND_657[184:0];
  _RAND_658 = {6{`RANDOM}};
  cache_data_655 = _RAND_658[184:0];
  _RAND_659 = {6{`RANDOM}};
  cache_data_656 = _RAND_659[184:0];
  _RAND_660 = {6{`RANDOM}};
  cache_data_657 = _RAND_660[184:0];
  _RAND_661 = {6{`RANDOM}};
  cache_data_658 = _RAND_661[184:0];
  _RAND_662 = {6{`RANDOM}};
  cache_data_659 = _RAND_662[184:0];
  _RAND_663 = {6{`RANDOM}};
  cache_data_660 = _RAND_663[184:0];
  _RAND_664 = {6{`RANDOM}};
  cache_data_661 = _RAND_664[184:0];
  _RAND_665 = {6{`RANDOM}};
  cache_data_662 = _RAND_665[184:0];
  _RAND_666 = {6{`RANDOM}};
  cache_data_663 = _RAND_666[184:0];
  _RAND_667 = {6{`RANDOM}};
  cache_data_664 = _RAND_667[184:0];
  _RAND_668 = {6{`RANDOM}};
  cache_data_665 = _RAND_668[184:0];
  _RAND_669 = {6{`RANDOM}};
  cache_data_666 = _RAND_669[184:0];
  _RAND_670 = {6{`RANDOM}};
  cache_data_667 = _RAND_670[184:0];
  _RAND_671 = {6{`RANDOM}};
  cache_data_668 = _RAND_671[184:0];
  _RAND_672 = {6{`RANDOM}};
  cache_data_669 = _RAND_672[184:0];
  _RAND_673 = {6{`RANDOM}};
  cache_data_670 = _RAND_673[184:0];
  _RAND_674 = {6{`RANDOM}};
  cache_data_671 = _RAND_674[184:0];
  _RAND_675 = {6{`RANDOM}};
  cache_data_672 = _RAND_675[184:0];
  _RAND_676 = {6{`RANDOM}};
  cache_data_673 = _RAND_676[184:0];
  _RAND_677 = {6{`RANDOM}};
  cache_data_674 = _RAND_677[184:0];
  _RAND_678 = {6{`RANDOM}};
  cache_data_675 = _RAND_678[184:0];
  _RAND_679 = {6{`RANDOM}};
  cache_data_676 = _RAND_679[184:0];
  _RAND_680 = {6{`RANDOM}};
  cache_data_677 = _RAND_680[184:0];
  _RAND_681 = {6{`RANDOM}};
  cache_data_678 = _RAND_681[184:0];
  _RAND_682 = {6{`RANDOM}};
  cache_data_679 = _RAND_682[184:0];
  _RAND_683 = {6{`RANDOM}};
  cache_data_680 = _RAND_683[184:0];
  _RAND_684 = {6{`RANDOM}};
  cache_data_681 = _RAND_684[184:0];
  _RAND_685 = {6{`RANDOM}};
  cache_data_682 = _RAND_685[184:0];
  _RAND_686 = {6{`RANDOM}};
  cache_data_683 = _RAND_686[184:0];
  _RAND_687 = {6{`RANDOM}};
  cache_data_684 = _RAND_687[184:0];
  _RAND_688 = {6{`RANDOM}};
  cache_data_685 = _RAND_688[184:0];
  _RAND_689 = {6{`RANDOM}};
  cache_data_686 = _RAND_689[184:0];
  _RAND_690 = {6{`RANDOM}};
  cache_data_687 = _RAND_690[184:0];
  _RAND_691 = {6{`RANDOM}};
  cache_data_688 = _RAND_691[184:0];
  _RAND_692 = {6{`RANDOM}};
  cache_data_689 = _RAND_692[184:0];
  _RAND_693 = {6{`RANDOM}};
  cache_data_690 = _RAND_693[184:0];
  _RAND_694 = {6{`RANDOM}};
  cache_data_691 = _RAND_694[184:0];
  _RAND_695 = {6{`RANDOM}};
  cache_data_692 = _RAND_695[184:0];
  _RAND_696 = {6{`RANDOM}};
  cache_data_693 = _RAND_696[184:0];
  _RAND_697 = {6{`RANDOM}};
  cache_data_694 = _RAND_697[184:0];
  _RAND_698 = {6{`RANDOM}};
  cache_data_695 = _RAND_698[184:0];
  _RAND_699 = {6{`RANDOM}};
  cache_data_696 = _RAND_699[184:0];
  _RAND_700 = {6{`RANDOM}};
  cache_data_697 = _RAND_700[184:0];
  _RAND_701 = {6{`RANDOM}};
  cache_data_698 = _RAND_701[184:0];
  _RAND_702 = {6{`RANDOM}};
  cache_data_699 = _RAND_702[184:0];
  _RAND_703 = {6{`RANDOM}};
  cache_data_700 = _RAND_703[184:0];
  _RAND_704 = {6{`RANDOM}};
  cache_data_701 = _RAND_704[184:0];
  _RAND_705 = {6{`RANDOM}};
  cache_data_702 = _RAND_705[184:0];
  _RAND_706 = {6{`RANDOM}};
  cache_data_703 = _RAND_706[184:0];
  _RAND_707 = {6{`RANDOM}};
  cache_data_704 = _RAND_707[184:0];
  _RAND_708 = {6{`RANDOM}};
  cache_data_705 = _RAND_708[184:0];
  _RAND_709 = {6{`RANDOM}};
  cache_data_706 = _RAND_709[184:0];
  _RAND_710 = {6{`RANDOM}};
  cache_data_707 = _RAND_710[184:0];
  _RAND_711 = {6{`RANDOM}};
  cache_data_708 = _RAND_711[184:0];
  _RAND_712 = {6{`RANDOM}};
  cache_data_709 = _RAND_712[184:0];
  _RAND_713 = {6{`RANDOM}};
  cache_data_710 = _RAND_713[184:0];
  _RAND_714 = {6{`RANDOM}};
  cache_data_711 = _RAND_714[184:0];
  _RAND_715 = {6{`RANDOM}};
  cache_data_712 = _RAND_715[184:0];
  _RAND_716 = {6{`RANDOM}};
  cache_data_713 = _RAND_716[184:0];
  _RAND_717 = {6{`RANDOM}};
  cache_data_714 = _RAND_717[184:0];
  _RAND_718 = {6{`RANDOM}};
  cache_data_715 = _RAND_718[184:0];
  _RAND_719 = {6{`RANDOM}};
  cache_data_716 = _RAND_719[184:0];
  _RAND_720 = {6{`RANDOM}};
  cache_data_717 = _RAND_720[184:0];
  _RAND_721 = {6{`RANDOM}};
  cache_data_718 = _RAND_721[184:0];
  _RAND_722 = {6{`RANDOM}};
  cache_data_719 = _RAND_722[184:0];
  _RAND_723 = {6{`RANDOM}};
  cache_data_720 = _RAND_723[184:0];
  _RAND_724 = {6{`RANDOM}};
  cache_data_721 = _RAND_724[184:0];
  _RAND_725 = {6{`RANDOM}};
  cache_data_722 = _RAND_725[184:0];
  _RAND_726 = {6{`RANDOM}};
  cache_data_723 = _RAND_726[184:0];
  _RAND_727 = {6{`RANDOM}};
  cache_data_724 = _RAND_727[184:0];
  _RAND_728 = {6{`RANDOM}};
  cache_data_725 = _RAND_728[184:0];
  _RAND_729 = {6{`RANDOM}};
  cache_data_726 = _RAND_729[184:0];
  _RAND_730 = {6{`RANDOM}};
  cache_data_727 = _RAND_730[184:0];
  _RAND_731 = {6{`RANDOM}};
  cache_data_728 = _RAND_731[184:0];
  _RAND_732 = {6{`RANDOM}};
  cache_data_729 = _RAND_732[184:0];
  _RAND_733 = {6{`RANDOM}};
  cache_data_730 = _RAND_733[184:0];
  _RAND_734 = {6{`RANDOM}};
  cache_data_731 = _RAND_734[184:0];
  _RAND_735 = {6{`RANDOM}};
  cache_data_732 = _RAND_735[184:0];
  _RAND_736 = {6{`RANDOM}};
  cache_data_733 = _RAND_736[184:0];
  _RAND_737 = {6{`RANDOM}};
  cache_data_734 = _RAND_737[184:0];
  _RAND_738 = {6{`RANDOM}};
  cache_data_735 = _RAND_738[184:0];
  _RAND_739 = {6{`RANDOM}};
  cache_data_736 = _RAND_739[184:0];
  _RAND_740 = {6{`RANDOM}};
  cache_data_737 = _RAND_740[184:0];
  _RAND_741 = {6{`RANDOM}};
  cache_data_738 = _RAND_741[184:0];
  _RAND_742 = {6{`RANDOM}};
  cache_data_739 = _RAND_742[184:0];
  _RAND_743 = {6{`RANDOM}};
  cache_data_740 = _RAND_743[184:0];
  _RAND_744 = {6{`RANDOM}};
  cache_data_741 = _RAND_744[184:0];
  _RAND_745 = {6{`RANDOM}};
  cache_data_742 = _RAND_745[184:0];
  _RAND_746 = {6{`RANDOM}};
  cache_data_743 = _RAND_746[184:0];
  _RAND_747 = {6{`RANDOM}};
  cache_data_744 = _RAND_747[184:0];
  _RAND_748 = {6{`RANDOM}};
  cache_data_745 = _RAND_748[184:0];
  _RAND_749 = {6{`RANDOM}};
  cache_data_746 = _RAND_749[184:0];
  _RAND_750 = {6{`RANDOM}};
  cache_data_747 = _RAND_750[184:0];
  _RAND_751 = {6{`RANDOM}};
  cache_data_748 = _RAND_751[184:0];
  _RAND_752 = {6{`RANDOM}};
  cache_data_749 = _RAND_752[184:0];
  _RAND_753 = {6{`RANDOM}};
  cache_data_750 = _RAND_753[184:0];
  _RAND_754 = {6{`RANDOM}};
  cache_data_751 = _RAND_754[184:0];
  _RAND_755 = {6{`RANDOM}};
  cache_data_752 = _RAND_755[184:0];
  _RAND_756 = {6{`RANDOM}};
  cache_data_753 = _RAND_756[184:0];
  _RAND_757 = {6{`RANDOM}};
  cache_data_754 = _RAND_757[184:0];
  _RAND_758 = {6{`RANDOM}};
  cache_data_755 = _RAND_758[184:0];
  _RAND_759 = {6{`RANDOM}};
  cache_data_756 = _RAND_759[184:0];
  _RAND_760 = {6{`RANDOM}};
  cache_data_757 = _RAND_760[184:0];
  _RAND_761 = {6{`RANDOM}};
  cache_data_758 = _RAND_761[184:0];
  _RAND_762 = {6{`RANDOM}};
  cache_data_759 = _RAND_762[184:0];
  _RAND_763 = {6{`RANDOM}};
  cache_data_760 = _RAND_763[184:0];
  _RAND_764 = {6{`RANDOM}};
  cache_data_761 = _RAND_764[184:0];
  _RAND_765 = {6{`RANDOM}};
  cache_data_762 = _RAND_765[184:0];
  _RAND_766 = {6{`RANDOM}};
  cache_data_763 = _RAND_766[184:0];
  _RAND_767 = {6{`RANDOM}};
  cache_data_764 = _RAND_767[184:0];
  _RAND_768 = {6{`RANDOM}};
  cache_data_765 = _RAND_768[184:0];
  _RAND_769 = {6{`RANDOM}};
  cache_data_766 = _RAND_769[184:0];
  _RAND_770 = {6{`RANDOM}};
  cache_data_767 = _RAND_770[184:0];
  _RAND_771 = {6{`RANDOM}};
  cache_data_768 = _RAND_771[184:0];
  _RAND_772 = {6{`RANDOM}};
  cache_data_769 = _RAND_772[184:0];
  _RAND_773 = {6{`RANDOM}};
  cache_data_770 = _RAND_773[184:0];
  _RAND_774 = {6{`RANDOM}};
  cache_data_771 = _RAND_774[184:0];
  _RAND_775 = {6{`RANDOM}};
  cache_data_772 = _RAND_775[184:0];
  _RAND_776 = {6{`RANDOM}};
  cache_data_773 = _RAND_776[184:0];
  _RAND_777 = {6{`RANDOM}};
  cache_data_774 = _RAND_777[184:0];
  _RAND_778 = {6{`RANDOM}};
  cache_data_775 = _RAND_778[184:0];
  _RAND_779 = {6{`RANDOM}};
  cache_data_776 = _RAND_779[184:0];
  _RAND_780 = {6{`RANDOM}};
  cache_data_777 = _RAND_780[184:0];
  _RAND_781 = {6{`RANDOM}};
  cache_data_778 = _RAND_781[184:0];
  _RAND_782 = {6{`RANDOM}};
  cache_data_779 = _RAND_782[184:0];
  _RAND_783 = {6{`RANDOM}};
  cache_data_780 = _RAND_783[184:0];
  _RAND_784 = {6{`RANDOM}};
  cache_data_781 = _RAND_784[184:0];
  _RAND_785 = {6{`RANDOM}};
  cache_data_782 = _RAND_785[184:0];
  _RAND_786 = {6{`RANDOM}};
  cache_data_783 = _RAND_786[184:0];
  _RAND_787 = {6{`RANDOM}};
  cache_data_784 = _RAND_787[184:0];
  _RAND_788 = {6{`RANDOM}};
  cache_data_785 = _RAND_788[184:0];
  _RAND_789 = {6{`RANDOM}};
  cache_data_786 = _RAND_789[184:0];
  _RAND_790 = {6{`RANDOM}};
  cache_data_787 = _RAND_790[184:0];
  _RAND_791 = {6{`RANDOM}};
  cache_data_788 = _RAND_791[184:0];
  _RAND_792 = {6{`RANDOM}};
  cache_data_789 = _RAND_792[184:0];
  _RAND_793 = {6{`RANDOM}};
  cache_data_790 = _RAND_793[184:0];
  _RAND_794 = {6{`RANDOM}};
  cache_data_791 = _RAND_794[184:0];
  _RAND_795 = {6{`RANDOM}};
  cache_data_792 = _RAND_795[184:0];
  _RAND_796 = {6{`RANDOM}};
  cache_data_793 = _RAND_796[184:0];
  _RAND_797 = {6{`RANDOM}};
  cache_data_794 = _RAND_797[184:0];
  _RAND_798 = {6{`RANDOM}};
  cache_data_795 = _RAND_798[184:0];
  _RAND_799 = {6{`RANDOM}};
  cache_data_796 = _RAND_799[184:0];
  _RAND_800 = {6{`RANDOM}};
  cache_data_797 = _RAND_800[184:0];
  _RAND_801 = {6{`RANDOM}};
  cache_data_798 = _RAND_801[184:0];
  _RAND_802 = {6{`RANDOM}};
  cache_data_799 = _RAND_802[184:0];
  _RAND_803 = {6{`RANDOM}};
  cache_data_800 = _RAND_803[184:0];
  _RAND_804 = {6{`RANDOM}};
  cache_data_801 = _RAND_804[184:0];
  _RAND_805 = {6{`RANDOM}};
  cache_data_802 = _RAND_805[184:0];
  _RAND_806 = {6{`RANDOM}};
  cache_data_803 = _RAND_806[184:0];
  _RAND_807 = {6{`RANDOM}};
  cache_data_804 = _RAND_807[184:0];
  _RAND_808 = {6{`RANDOM}};
  cache_data_805 = _RAND_808[184:0];
  _RAND_809 = {6{`RANDOM}};
  cache_data_806 = _RAND_809[184:0];
  _RAND_810 = {6{`RANDOM}};
  cache_data_807 = _RAND_810[184:0];
  _RAND_811 = {6{`RANDOM}};
  cache_data_808 = _RAND_811[184:0];
  _RAND_812 = {6{`RANDOM}};
  cache_data_809 = _RAND_812[184:0];
  _RAND_813 = {6{`RANDOM}};
  cache_data_810 = _RAND_813[184:0];
  _RAND_814 = {6{`RANDOM}};
  cache_data_811 = _RAND_814[184:0];
  _RAND_815 = {6{`RANDOM}};
  cache_data_812 = _RAND_815[184:0];
  _RAND_816 = {6{`RANDOM}};
  cache_data_813 = _RAND_816[184:0];
  _RAND_817 = {6{`RANDOM}};
  cache_data_814 = _RAND_817[184:0];
  _RAND_818 = {6{`RANDOM}};
  cache_data_815 = _RAND_818[184:0];
  _RAND_819 = {6{`RANDOM}};
  cache_data_816 = _RAND_819[184:0];
  _RAND_820 = {6{`RANDOM}};
  cache_data_817 = _RAND_820[184:0];
  _RAND_821 = {6{`RANDOM}};
  cache_data_818 = _RAND_821[184:0];
  _RAND_822 = {6{`RANDOM}};
  cache_data_819 = _RAND_822[184:0];
  _RAND_823 = {6{`RANDOM}};
  cache_data_820 = _RAND_823[184:0];
  _RAND_824 = {6{`RANDOM}};
  cache_data_821 = _RAND_824[184:0];
  _RAND_825 = {6{`RANDOM}};
  cache_data_822 = _RAND_825[184:0];
  _RAND_826 = {6{`RANDOM}};
  cache_data_823 = _RAND_826[184:0];
  _RAND_827 = {6{`RANDOM}};
  cache_data_824 = _RAND_827[184:0];
  _RAND_828 = {6{`RANDOM}};
  cache_data_825 = _RAND_828[184:0];
  _RAND_829 = {6{`RANDOM}};
  cache_data_826 = _RAND_829[184:0];
  _RAND_830 = {6{`RANDOM}};
  cache_data_827 = _RAND_830[184:0];
  _RAND_831 = {6{`RANDOM}};
  cache_data_828 = _RAND_831[184:0];
  _RAND_832 = {6{`RANDOM}};
  cache_data_829 = _RAND_832[184:0];
  _RAND_833 = {6{`RANDOM}};
  cache_data_830 = _RAND_833[184:0];
  _RAND_834 = {6{`RANDOM}};
  cache_data_831 = _RAND_834[184:0];
  _RAND_835 = {6{`RANDOM}};
  cache_data_832 = _RAND_835[184:0];
  _RAND_836 = {6{`RANDOM}};
  cache_data_833 = _RAND_836[184:0];
  _RAND_837 = {6{`RANDOM}};
  cache_data_834 = _RAND_837[184:0];
  _RAND_838 = {6{`RANDOM}};
  cache_data_835 = _RAND_838[184:0];
  _RAND_839 = {6{`RANDOM}};
  cache_data_836 = _RAND_839[184:0];
  _RAND_840 = {6{`RANDOM}};
  cache_data_837 = _RAND_840[184:0];
  _RAND_841 = {6{`RANDOM}};
  cache_data_838 = _RAND_841[184:0];
  _RAND_842 = {6{`RANDOM}};
  cache_data_839 = _RAND_842[184:0];
  _RAND_843 = {6{`RANDOM}};
  cache_data_840 = _RAND_843[184:0];
  _RAND_844 = {6{`RANDOM}};
  cache_data_841 = _RAND_844[184:0];
  _RAND_845 = {6{`RANDOM}};
  cache_data_842 = _RAND_845[184:0];
  _RAND_846 = {6{`RANDOM}};
  cache_data_843 = _RAND_846[184:0];
  _RAND_847 = {6{`RANDOM}};
  cache_data_844 = _RAND_847[184:0];
  _RAND_848 = {6{`RANDOM}};
  cache_data_845 = _RAND_848[184:0];
  _RAND_849 = {6{`RANDOM}};
  cache_data_846 = _RAND_849[184:0];
  _RAND_850 = {6{`RANDOM}};
  cache_data_847 = _RAND_850[184:0];
  _RAND_851 = {6{`RANDOM}};
  cache_data_848 = _RAND_851[184:0];
  _RAND_852 = {6{`RANDOM}};
  cache_data_849 = _RAND_852[184:0];
  _RAND_853 = {6{`RANDOM}};
  cache_data_850 = _RAND_853[184:0];
  _RAND_854 = {6{`RANDOM}};
  cache_data_851 = _RAND_854[184:0];
  _RAND_855 = {6{`RANDOM}};
  cache_data_852 = _RAND_855[184:0];
  _RAND_856 = {6{`RANDOM}};
  cache_data_853 = _RAND_856[184:0];
  _RAND_857 = {6{`RANDOM}};
  cache_data_854 = _RAND_857[184:0];
  _RAND_858 = {6{`RANDOM}};
  cache_data_855 = _RAND_858[184:0];
  _RAND_859 = {6{`RANDOM}};
  cache_data_856 = _RAND_859[184:0];
  _RAND_860 = {6{`RANDOM}};
  cache_data_857 = _RAND_860[184:0];
  _RAND_861 = {6{`RANDOM}};
  cache_data_858 = _RAND_861[184:0];
  _RAND_862 = {6{`RANDOM}};
  cache_data_859 = _RAND_862[184:0];
  _RAND_863 = {6{`RANDOM}};
  cache_data_860 = _RAND_863[184:0];
  _RAND_864 = {6{`RANDOM}};
  cache_data_861 = _RAND_864[184:0];
  _RAND_865 = {6{`RANDOM}};
  cache_data_862 = _RAND_865[184:0];
  _RAND_866 = {6{`RANDOM}};
  cache_data_863 = _RAND_866[184:0];
  _RAND_867 = {6{`RANDOM}};
  cache_data_864 = _RAND_867[184:0];
  _RAND_868 = {6{`RANDOM}};
  cache_data_865 = _RAND_868[184:0];
  _RAND_869 = {6{`RANDOM}};
  cache_data_866 = _RAND_869[184:0];
  _RAND_870 = {6{`RANDOM}};
  cache_data_867 = _RAND_870[184:0];
  _RAND_871 = {6{`RANDOM}};
  cache_data_868 = _RAND_871[184:0];
  _RAND_872 = {6{`RANDOM}};
  cache_data_869 = _RAND_872[184:0];
  _RAND_873 = {6{`RANDOM}};
  cache_data_870 = _RAND_873[184:0];
  _RAND_874 = {6{`RANDOM}};
  cache_data_871 = _RAND_874[184:0];
  _RAND_875 = {6{`RANDOM}};
  cache_data_872 = _RAND_875[184:0];
  _RAND_876 = {6{`RANDOM}};
  cache_data_873 = _RAND_876[184:0];
  _RAND_877 = {6{`RANDOM}};
  cache_data_874 = _RAND_877[184:0];
  _RAND_878 = {6{`RANDOM}};
  cache_data_875 = _RAND_878[184:0];
  _RAND_879 = {6{`RANDOM}};
  cache_data_876 = _RAND_879[184:0];
  _RAND_880 = {6{`RANDOM}};
  cache_data_877 = _RAND_880[184:0];
  _RAND_881 = {6{`RANDOM}};
  cache_data_878 = _RAND_881[184:0];
  _RAND_882 = {6{`RANDOM}};
  cache_data_879 = _RAND_882[184:0];
  _RAND_883 = {6{`RANDOM}};
  cache_data_880 = _RAND_883[184:0];
  _RAND_884 = {6{`RANDOM}};
  cache_data_881 = _RAND_884[184:0];
  _RAND_885 = {6{`RANDOM}};
  cache_data_882 = _RAND_885[184:0];
  _RAND_886 = {6{`RANDOM}};
  cache_data_883 = _RAND_886[184:0];
  _RAND_887 = {6{`RANDOM}};
  cache_data_884 = _RAND_887[184:0];
  _RAND_888 = {6{`RANDOM}};
  cache_data_885 = _RAND_888[184:0];
  _RAND_889 = {6{`RANDOM}};
  cache_data_886 = _RAND_889[184:0];
  _RAND_890 = {6{`RANDOM}};
  cache_data_887 = _RAND_890[184:0];
  _RAND_891 = {6{`RANDOM}};
  cache_data_888 = _RAND_891[184:0];
  _RAND_892 = {6{`RANDOM}};
  cache_data_889 = _RAND_892[184:0];
  _RAND_893 = {6{`RANDOM}};
  cache_data_890 = _RAND_893[184:0];
  _RAND_894 = {6{`RANDOM}};
  cache_data_891 = _RAND_894[184:0];
  _RAND_895 = {6{`RANDOM}};
  cache_data_892 = _RAND_895[184:0];
  _RAND_896 = {6{`RANDOM}};
  cache_data_893 = _RAND_896[184:0];
  _RAND_897 = {6{`RANDOM}};
  cache_data_894 = _RAND_897[184:0];
  _RAND_898 = {6{`RANDOM}};
  cache_data_895 = _RAND_898[184:0];
  _RAND_899 = {6{`RANDOM}};
  cache_data_896 = _RAND_899[184:0];
  _RAND_900 = {6{`RANDOM}};
  cache_data_897 = _RAND_900[184:0];
  _RAND_901 = {6{`RANDOM}};
  cache_data_898 = _RAND_901[184:0];
  _RAND_902 = {6{`RANDOM}};
  cache_data_899 = _RAND_902[184:0];
  _RAND_903 = {6{`RANDOM}};
  cache_data_900 = _RAND_903[184:0];
  _RAND_904 = {6{`RANDOM}};
  cache_data_901 = _RAND_904[184:0];
  _RAND_905 = {6{`RANDOM}};
  cache_data_902 = _RAND_905[184:0];
  _RAND_906 = {6{`RANDOM}};
  cache_data_903 = _RAND_906[184:0];
  _RAND_907 = {6{`RANDOM}};
  cache_data_904 = _RAND_907[184:0];
  _RAND_908 = {6{`RANDOM}};
  cache_data_905 = _RAND_908[184:0];
  _RAND_909 = {6{`RANDOM}};
  cache_data_906 = _RAND_909[184:0];
  _RAND_910 = {6{`RANDOM}};
  cache_data_907 = _RAND_910[184:0];
  _RAND_911 = {6{`RANDOM}};
  cache_data_908 = _RAND_911[184:0];
  _RAND_912 = {6{`RANDOM}};
  cache_data_909 = _RAND_912[184:0];
  _RAND_913 = {6{`RANDOM}};
  cache_data_910 = _RAND_913[184:0];
  _RAND_914 = {6{`RANDOM}};
  cache_data_911 = _RAND_914[184:0];
  _RAND_915 = {6{`RANDOM}};
  cache_data_912 = _RAND_915[184:0];
  _RAND_916 = {6{`RANDOM}};
  cache_data_913 = _RAND_916[184:0];
  _RAND_917 = {6{`RANDOM}};
  cache_data_914 = _RAND_917[184:0];
  _RAND_918 = {6{`RANDOM}};
  cache_data_915 = _RAND_918[184:0];
  _RAND_919 = {6{`RANDOM}};
  cache_data_916 = _RAND_919[184:0];
  _RAND_920 = {6{`RANDOM}};
  cache_data_917 = _RAND_920[184:0];
  _RAND_921 = {6{`RANDOM}};
  cache_data_918 = _RAND_921[184:0];
  _RAND_922 = {6{`RANDOM}};
  cache_data_919 = _RAND_922[184:0];
  _RAND_923 = {6{`RANDOM}};
  cache_data_920 = _RAND_923[184:0];
  _RAND_924 = {6{`RANDOM}};
  cache_data_921 = _RAND_924[184:0];
  _RAND_925 = {6{`RANDOM}};
  cache_data_922 = _RAND_925[184:0];
  _RAND_926 = {6{`RANDOM}};
  cache_data_923 = _RAND_926[184:0];
  _RAND_927 = {6{`RANDOM}};
  cache_data_924 = _RAND_927[184:0];
  _RAND_928 = {6{`RANDOM}};
  cache_data_925 = _RAND_928[184:0];
  _RAND_929 = {6{`RANDOM}};
  cache_data_926 = _RAND_929[184:0];
  _RAND_930 = {6{`RANDOM}};
  cache_data_927 = _RAND_930[184:0];
  _RAND_931 = {6{`RANDOM}};
  cache_data_928 = _RAND_931[184:0];
  _RAND_932 = {6{`RANDOM}};
  cache_data_929 = _RAND_932[184:0];
  _RAND_933 = {6{`RANDOM}};
  cache_data_930 = _RAND_933[184:0];
  _RAND_934 = {6{`RANDOM}};
  cache_data_931 = _RAND_934[184:0];
  _RAND_935 = {6{`RANDOM}};
  cache_data_932 = _RAND_935[184:0];
  _RAND_936 = {6{`RANDOM}};
  cache_data_933 = _RAND_936[184:0];
  _RAND_937 = {6{`RANDOM}};
  cache_data_934 = _RAND_937[184:0];
  _RAND_938 = {6{`RANDOM}};
  cache_data_935 = _RAND_938[184:0];
  _RAND_939 = {6{`RANDOM}};
  cache_data_936 = _RAND_939[184:0];
  _RAND_940 = {6{`RANDOM}};
  cache_data_937 = _RAND_940[184:0];
  _RAND_941 = {6{`RANDOM}};
  cache_data_938 = _RAND_941[184:0];
  _RAND_942 = {6{`RANDOM}};
  cache_data_939 = _RAND_942[184:0];
  _RAND_943 = {6{`RANDOM}};
  cache_data_940 = _RAND_943[184:0];
  _RAND_944 = {6{`RANDOM}};
  cache_data_941 = _RAND_944[184:0];
  _RAND_945 = {6{`RANDOM}};
  cache_data_942 = _RAND_945[184:0];
  _RAND_946 = {6{`RANDOM}};
  cache_data_943 = _RAND_946[184:0];
  _RAND_947 = {6{`RANDOM}};
  cache_data_944 = _RAND_947[184:0];
  _RAND_948 = {6{`RANDOM}};
  cache_data_945 = _RAND_948[184:0];
  _RAND_949 = {6{`RANDOM}};
  cache_data_946 = _RAND_949[184:0];
  _RAND_950 = {6{`RANDOM}};
  cache_data_947 = _RAND_950[184:0];
  _RAND_951 = {6{`RANDOM}};
  cache_data_948 = _RAND_951[184:0];
  _RAND_952 = {6{`RANDOM}};
  cache_data_949 = _RAND_952[184:0];
  _RAND_953 = {6{`RANDOM}};
  cache_data_950 = _RAND_953[184:0];
  _RAND_954 = {6{`RANDOM}};
  cache_data_951 = _RAND_954[184:0];
  _RAND_955 = {6{`RANDOM}};
  cache_data_952 = _RAND_955[184:0];
  _RAND_956 = {6{`RANDOM}};
  cache_data_953 = _RAND_956[184:0];
  _RAND_957 = {6{`RANDOM}};
  cache_data_954 = _RAND_957[184:0];
  _RAND_958 = {6{`RANDOM}};
  cache_data_955 = _RAND_958[184:0];
  _RAND_959 = {6{`RANDOM}};
  cache_data_956 = _RAND_959[184:0];
  _RAND_960 = {6{`RANDOM}};
  cache_data_957 = _RAND_960[184:0];
  _RAND_961 = {6{`RANDOM}};
  cache_data_958 = _RAND_961[184:0];
  _RAND_962 = {6{`RANDOM}};
  cache_data_959 = _RAND_962[184:0];
  _RAND_963 = {6{`RANDOM}};
  cache_data_960 = _RAND_963[184:0];
  _RAND_964 = {6{`RANDOM}};
  cache_data_961 = _RAND_964[184:0];
  _RAND_965 = {6{`RANDOM}};
  cache_data_962 = _RAND_965[184:0];
  _RAND_966 = {6{`RANDOM}};
  cache_data_963 = _RAND_966[184:0];
  _RAND_967 = {6{`RANDOM}};
  cache_data_964 = _RAND_967[184:0];
  _RAND_968 = {6{`RANDOM}};
  cache_data_965 = _RAND_968[184:0];
  _RAND_969 = {6{`RANDOM}};
  cache_data_966 = _RAND_969[184:0];
  _RAND_970 = {6{`RANDOM}};
  cache_data_967 = _RAND_970[184:0];
  _RAND_971 = {6{`RANDOM}};
  cache_data_968 = _RAND_971[184:0];
  _RAND_972 = {6{`RANDOM}};
  cache_data_969 = _RAND_972[184:0];
  _RAND_973 = {6{`RANDOM}};
  cache_data_970 = _RAND_973[184:0];
  _RAND_974 = {6{`RANDOM}};
  cache_data_971 = _RAND_974[184:0];
  _RAND_975 = {6{`RANDOM}};
  cache_data_972 = _RAND_975[184:0];
  _RAND_976 = {6{`RANDOM}};
  cache_data_973 = _RAND_976[184:0];
  _RAND_977 = {6{`RANDOM}};
  cache_data_974 = _RAND_977[184:0];
  _RAND_978 = {6{`RANDOM}};
  cache_data_975 = _RAND_978[184:0];
  _RAND_979 = {6{`RANDOM}};
  cache_data_976 = _RAND_979[184:0];
  _RAND_980 = {6{`RANDOM}};
  cache_data_977 = _RAND_980[184:0];
  _RAND_981 = {6{`RANDOM}};
  cache_data_978 = _RAND_981[184:0];
  _RAND_982 = {6{`RANDOM}};
  cache_data_979 = _RAND_982[184:0];
  _RAND_983 = {6{`RANDOM}};
  cache_data_980 = _RAND_983[184:0];
  _RAND_984 = {6{`RANDOM}};
  cache_data_981 = _RAND_984[184:0];
  _RAND_985 = {6{`RANDOM}};
  cache_data_982 = _RAND_985[184:0];
  _RAND_986 = {6{`RANDOM}};
  cache_data_983 = _RAND_986[184:0];
  _RAND_987 = {6{`RANDOM}};
  cache_data_984 = _RAND_987[184:0];
  _RAND_988 = {6{`RANDOM}};
  cache_data_985 = _RAND_988[184:0];
  _RAND_989 = {6{`RANDOM}};
  cache_data_986 = _RAND_989[184:0];
  _RAND_990 = {6{`RANDOM}};
  cache_data_987 = _RAND_990[184:0];
  _RAND_991 = {6{`RANDOM}};
  cache_data_988 = _RAND_991[184:0];
  _RAND_992 = {6{`RANDOM}};
  cache_data_989 = _RAND_992[184:0];
  _RAND_993 = {6{`RANDOM}};
  cache_data_990 = _RAND_993[184:0];
  _RAND_994 = {6{`RANDOM}};
  cache_data_991 = _RAND_994[184:0];
  _RAND_995 = {6{`RANDOM}};
  cache_data_992 = _RAND_995[184:0];
  _RAND_996 = {6{`RANDOM}};
  cache_data_993 = _RAND_996[184:0];
  _RAND_997 = {6{`RANDOM}};
  cache_data_994 = _RAND_997[184:0];
  _RAND_998 = {6{`RANDOM}};
  cache_data_995 = _RAND_998[184:0];
  _RAND_999 = {6{`RANDOM}};
  cache_data_996 = _RAND_999[184:0];
  _RAND_1000 = {6{`RANDOM}};
  cache_data_997 = _RAND_1000[184:0];
  _RAND_1001 = {6{`RANDOM}};
  cache_data_998 = _RAND_1001[184:0];
  _RAND_1002 = {6{`RANDOM}};
  cache_data_999 = _RAND_1002[184:0];
  _RAND_1003 = {6{`RANDOM}};
  cache_data_1000 = _RAND_1003[184:0];
  _RAND_1004 = {6{`RANDOM}};
  cache_data_1001 = _RAND_1004[184:0];
  _RAND_1005 = {6{`RANDOM}};
  cache_data_1002 = _RAND_1005[184:0];
  _RAND_1006 = {6{`RANDOM}};
  cache_data_1003 = _RAND_1006[184:0];
  _RAND_1007 = {6{`RANDOM}};
  cache_data_1004 = _RAND_1007[184:0];
  _RAND_1008 = {6{`RANDOM}};
  cache_data_1005 = _RAND_1008[184:0];
  _RAND_1009 = {6{`RANDOM}};
  cache_data_1006 = _RAND_1009[184:0];
  _RAND_1010 = {6{`RANDOM}};
  cache_data_1007 = _RAND_1010[184:0];
  _RAND_1011 = {6{`RANDOM}};
  cache_data_1008 = _RAND_1011[184:0];
  _RAND_1012 = {6{`RANDOM}};
  cache_data_1009 = _RAND_1012[184:0];
  _RAND_1013 = {6{`RANDOM}};
  cache_data_1010 = _RAND_1013[184:0];
  _RAND_1014 = {6{`RANDOM}};
  cache_data_1011 = _RAND_1014[184:0];
  _RAND_1015 = {6{`RANDOM}};
  cache_data_1012 = _RAND_1015[184:0];
  _RAND_1016 = {6{`RANDOM}};
  cache_data_1013 = _RAND_1016[184:0];
  _RAND_1017 = {6{`RANDOM}};
  cache_data_1014 = _RAND_1017[184:0];
  _RAND_1018 = {6{`RANDOM}};
  cache_data_1015 = _RAND_1018[184:0];
  _RAND_1019 = {6{`RANDOM}};
  cache_data_1016 = _RAND_1019[184:0];
  _RAND_1020 = {6{`RANDOM}};
  cache_data_1017 = _RAND_1020[184:0];
  _RAND_1021 = {6{`RANDOM}};
  cache_data_1018 = _RAND_1021[184:0];
  _RAND_1022 = {6{`RANDOM}};
  cache_data_1019 = _RAND_1022[184:0];
  _RAND_1023 = {6{`RANDOM}};
  cache_data_1020 = _RAND_1023[184:0];
  _RAND_1024 = {6{`RANDOM}};
  cache_data_1021 = _RAND_1024[184:0];
  _RAND_1025 = {6{`RANDOM}};
  cache_data_1022 = _RAND_1025[184:0];
  _RAND_1026 = {6{`RANDOM}};
  cache_data_1023 = _RAND_1026[184:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input         clock,
  input         reset,
  output [31:0] io_fs_pc,
  output [6:0]  io_op,
  output        io_in_WB,
  output [31:0] io_wb_pc,
  output [31:0] io_wb_inst,
  output [31:0] io_ds_pc,
  output [63:0] io_mem_result,
  output [2:0]  io_ld_type
);
  wire  ifu_clock; // @[TopMain.scala 23:23]
  wire  ifu_reset; // @[TopMain.scala 23:23]
  wire  ifu_io_reset; // @[TopMain.scala 23:23]
  wire [31:0] ifu_io_fd_bus_inst; // @[TopMain.scala 23:23]
  wire [31:0] ifu_io_fd_bus_pc; // @[TopMain.scala 23:23]
  wire  ifu_io_ds_allowin; // @[TopMain.scala 23:23]
  wire  ifu_io_fs_to_ds_valid; // @[TopMain.scala 23:23]
  wire  ifu_io_br_bus_br_taken; // @[TopMain.scala 23:23]
  wire [31:0] ifu_io_br_bus_br_target; // @[TopMain.scala 23:23]
  wire  ifu_io_br_bus_rawblock; // @[TopMain.scala 23:23]
  wire [63:0] ifu_io_br_bus_csr_rdata; // @[TopMain.scala 23:23]
  wire  ifu_io_br_bus_eval; // @[TopMain.scala 23:23]
  wire  ifu_io_br_bus_mret; // @[TopMain.scala 23:23]
  wire  ifu_io_inst_sram_req; // @[TopMain.scala 23:23]
  wire [63:0] ifu_io_inst_sram_addr; // @[TopMain.scala 23:23]
  wire [63:0] ifu_io_inst_sram_rdata; // @[TopMain.scala 23:23]
  wire  ifu_io_inst_sram_addr_ok; // @[TopMain.scala 23:23]
  wire  ifu_io_inst_sram_data_ok; // @[TopMain.scala 23:23]
  wire  idu_clock; // @[TopMain.scala 24:23]
  wire  idu_reset; // @[TopMain.scala 24:23]
  wire  idu_io_es_allowin; // @[TopMain.scala 24:23]
  wire  idu_io_ds_allowin; // @[TopMain.scala 24:23]
  wire  idu_io_fs_to_ds_valid; // @[TopMain.scala 24:23]
  wire  idu_io_ds_to_es_valid; // @[TopMain.scala 24:23]
  wire [31:0] idu_io_fd_bus_inst; // @[TopMain.scala 24:23]
  wire [31:0] idu_io_fd_bus_pc; // @[TopMain.scala 24:23]
  wire [7:0] idu_io_de_bus_OP; // @[TopMain.scala 24:23]
  wire  idu_io_de_bus_res_from_mem; // @[TopMain.scala 24:23]
  wire  idu_io_de_bus_gr_we; // @[TopMain.scala 24:23]
  wire  idu_io_de_bus_MemWen; // @[TopMain.scala 24:23]
  wire [7:0] idu_io_de_bus_wmask; // @[TopMain.scala 24:23]
  wire [31:0] idu_io_de_bus_ds_pc; // @[TopMain.scala 24:23]
  wire [4:0] idu_io_de_bus_dest; // @[TopMain.scala 24:23]
  wire [63:0] idu_io_de_bus_imm; // @[TopMain.scala 24:23]
  wire [63:0] idu_io_de_bus_rdata1; // @[TopMain.scala 24:23]
  wire [63:0] idu_io_de_bus_rdata2; // @[TopMain.scala 24:23]
  wire [2:0] idu_io_de_bus_ld_type; // @[TopMain.scala 24:23]
  wire [31:0] idu_io_de_bus_inst; // @[TopMain.scala 24:23]
  wire [63:0] idu_io_de_bus_csr_rdata; // @[TopMain.scala 24:23]
  wire [2:0] idu_io_de_bus_csr_waddr1; // @[TopMain.scala 24:23]
  wire [2:0] idu_io_de_bus_csr_waddr2; // @[TopMain.scala 24:23]
  wire [2:0] idu_io_de_bus_csr_raddr; // @[TopMain.scala 24:23]
  wire  idu_io_de_bus_csr_ren; // @[TopMain.scala 24:23]
  wire  idu_io_de_bus_csr_wen; // @[TopMain.scala 24:23]
  wire  idu_io_de_bus_eval; // @[TopMain.scala 24:23]
  wire  idu_io_de_bus_is_ld; // @[TopMain.scala 24:23]
  wire  idu_io_br_bus_br_taken; // @[TopMain.scala 24:23]
  wire [31:0] idu_io_br_bus_br_target; // @[TopMain.scala 24:23]
  wire  idu_io_br_bus_rawblock; // @[TopMain.scala 24:23]
  wire [63:0] idu_io_br_bus_csr_rdata; // @[TopMain.scala 24:23]
  wire  idu_io_br_bus_eval; // @[TopMain.scala 24:23]
  wire  idu_io_br_bus_mret; // @[TopMain.scala 24:23]
  wire  idu_io_rf_bus_rf_we; // @[TopMain.scala 24:23]
  wire [4:0] idu_io_rf_bus_rf_waddr; // @[TopMain.scala 24:23]
  wire [63:0] idu_io_rf_bus_rf_wdata; // @[TopMain.scala 24:23]
  wire [31:0] idu_io_rf_bus_wb_pc; // @[TopMain.scala 24:23]
  wire [31:0] idu_io_rf_bus_wb_inst; // @[TopMain.scala 24:23]
  wire [63:0] idu_io_rf_bus_csr_wdata; // @[TopMain.scala 24:23]
  wire  idu_io_rf_bus_csr_wen; // @[TopMain.scala 24:23]
  wire [2:0] idu_io_rf_bus_csr_waddr1; // @[TopMain.scala 24:23]
  wire [2:0] idu_io_rf_bus_csr_waddr2; // @[TopMain.scala 24:23]
  wire  idu_io_rf_bus_eval; // @[TopMain.scala 24:23]
  wire  idu_io_es_dest_valid_gr_we; // @[TopMain.scala 24:23]
  wire  idu_io_es_dest_valid_es_valid; // @[TopMain.scala 24:23]
  wire [4:0] idu_io_es_dest_valid_dest; // @[TopMain.scala 24:23]
  wire [63:0] idu_io_es_dest_valid_es_forward_data; // @[TopMain.scala 24:23]
  wire  idu_io_es_dest_valid_es_is_ld; // @[TopMain.scala 24:23]
  wire  idu_io_es_dest_valid_es_ready_go; // @[TopMain.scala 24:23]
  wire  idu_io_es_dest_valid_es_to_ms_valid; // @[TopMain.scala 24:23]
  wire  idu_io_ms_dest_valid_gr_we; // @[TopMain.scala 24:23]
  wire  idu_io_ms_dest_valid_ms_valid; // @[TopMain.scala 24:23]
  wire [4:0] idu_io_ms_dest_valid_dest; // @[TopMain.scala 24:23]
  wire [63:0] idu_io_ms_dest_valid_ms_forward_data; // @[TopMain.scala 24:23]
  wire  idu_io_ms_dest_valid_ms_is_ld; // @[TopMain.scala 24:23]
  wire  idu_io_ms_dest_valid_ms_to_ws_valid; // @[TopMain.scala 24:23]
  wire  idu_io_ms_dest_valid_ms_ready_go; // @[TopMain.scala 24:23]
  wire  idu_io_ws_dest_valid_gr_we; // @[TopMain.scala 24:23]
  wire  idu_io_ws_dest_valid_ws_valid; // @[TopMain.scala 24:23]
  wire [4:0] idu_io_ws_dest_valid_dest; // @[TopMain.scala 24:23]
  wire [63:0] idu_io_ws_dest_valid_ws_forward_data; // @[TopMain.scala 24:23]
  wire  exu_clock; // @[TopMain.scala 25:23]
  wire  exu_reset; // @[TopMain.scala 25:23]
  wire  exu_io_ms_allowin; // @[TopMain.scala 25:23]
  wire  exu_io_es_allowin; // @[TopMain.scala 25:23]
  wire  exu_io_ds_to_es_valid; // @[TopMain.scala 25:23]
  wire  exu_io_es_to_ms_valid; // @[TopMain.scala 25:23]
  wire [7:0] exu_io_de_bus_OP; // @[TopMain.scala 25:23]
  wire  exu_io_de_bus_res_from_mem; // @[TopMain.scala 25:23]
  wire  exu_io_de_bus_gr_we; // @[TopMain.scala 25:23]
  wire  exu_io_de_bus_MemWen; // @[TopMain.scala 25:23]
  wire [7:0] exu_io_de_bus_wmask; // @[TopMain.scala 25:23]
  wire [31:0] exu_io_de_bus_ds_pc; // @[TopMain.scala 25:23]
  wire [4:0] exu_io_de_bus_dest; // @[TopMain.scala 25:23]
  wire [63:0] exu_io_de_bus_imm; // @[TopMain.scala 25:23]
  wire [63:0] exu_io_de_bus_rdata1; // @[TopMain.scala 25:23]
  wire [63:0] exu_io_de_bus_rdata2; // @[TopMain.scala 25:23]
  wire [2:0] exu_io_de_bus_ld_type; // @[TopMain.scala 25:23]
  wire [31:0] exu_io_de_bus_inst; // @[TopMain.scala 25:23]
  wire [63:0] exu_io_de_bus_csr_rdata; // @[TopMain.scala 25:23]
  wire [2:0] exu_io_de_bus_csr_waddr1; // @[TopMain.scala 25:23]
  wire [2:0] exu_io_de_bus_csr_waddr2; // @[TopMain.scala 25:23]
  wire  exu_io_de_bus_csr_wen; // @[TopMain.scala 25:23]
  wire  exu_io_de_bus_eval; // @[TopMain.scala 25:23]
  wire  exu_io_de_bus_is_ld; // @[TopMain.scala 25:23]
  wire  exu_io_em_bus_res_from_mem; // @[TopMain.scala 25:23]
  wire  exu_io_em_bus_gr_we; // @[TopMain.scala 25:23]
  wire [4:0] exu_io_em_bus_dest; // @[TopMain.scala 25:23]
  wire [63:0] exu_io_em_bus_alu_result; // @[TopMain.scala 25:23]
  wire [31:0] exu_io_em_bus_ex_pc; // @[TopMain.scala 25:23]
  wire [2:0] exu_io_em_bus_ld_type; // @[TopMain.scala 25:23]
  wire [31:0] exu_io_em_bus_inst; // @[TopMain.scala 25:23]
  wire [63:0] exu_io_em_bus_csr_wdata; // @[TopMain.scala 25:23]
  wire  exu_io_em_bus_csr_wen; // @[TopMain.scala 25:23]
  wire [2:0] exu_io_em_bus_csr_waddr1; // @[TopMain.scala 25:23]
  wire [2:0] exu_io_em_bus_csr_waddr2; // @[TopMain.scala 25:23]
  wire  exu_io_em_bus_eval; // @[TopMain.scala 25:23]
  wire  exu_io_em_bus_is_ld; // @[TopMain.scala 25:23]
  wire  exu_io_em_bus_MemWen; // @[TopMain.scala 25:23]
  wire [63:0] exu_io_em_bus_Memwdata; // @[TopMain.scala 25:23]
  wire [7:0] exu_io_em_bus_wmask; // @[TopMain.scala 25:23]
  wire  exu_io_es_dest_valid_gr_we; // @[TopMain.scala 25:23]
  wire  exu_io_es_dest_valid_es_valid; // @[TopMain.scala 25:23]
  wire [4:0] exu_io_es_dest_valid_dest; // @[TopMain.scala 25:23]
  wire [63:0] exu_io_es_dest_valid_es_forward_data; // @[TopMain.scala 25:23]
  wire  exu_io_es_dest_valid_es_is_ld; // @[TopMain.scala 25:23]
  wire  exu_io_es_dest_valid_es_ready_go; // @[TopMain.scala 25:23]
  wire  exu_io_es_dest_valid_es_to_ms_valid; // @[TopMain.scala 25:23]
  wire  mem_clock; // @[TopMain.scala 26:23]
  wire  mem_reset; // @[TopMain.scala 26:23]
  wire  mem_io_ms_allowin; // @[TopMain.scala 26:23]
  wire  mem_io_es_to_ms_valid; // @[TopMain.scala 26:23]
  wire  mem_io_ms_to_ws_valid; // @[TopMain.scala 26:23]
  wire  mem_io_em_bus_res_from_mem; // @[TopMain.scala 26:23]
  wire  mem_io_em_bus_gr_we; // @[TopMain.scala 26:23]
  wire [4:0] mem_io_em_bus_dest; // @[TopMain.scala 26:23]
  wire [63:0] mem_io_em_bus_alu_result; // @[TopMain.scala 26:23]
  wire [31:0] mem_io_em_bus_ex_pc; // @[TopMain.scala 26:23]
  wire [2:0] mem_io_em_bus_ld_type; // @[TopMain.scala 26:23]
  wire [31:0] mem_io_em_bus_inst; // @[TopMain.scala 26:23]
  wire [63:0] mem_io_em_bus_csr_wdata; // @[TopMain.scala 26:23]
  wire  mem_io_em_bus_csr_wen; // @[TopMain.scala 26:23]
  wire [2:0] mem_io_em_bus_csr_waddr1; // @[TopMain.scala 26:23]
  wire [2:0] mem_io_em_bus_csr_waddr2; // @[TopMain.scala 26:23]
  wire  mem_io_em_bus_eval; // @[TopMain.scala 26:23]
  wire  mem_io_em_bus_is_ld; // @[TopMain.scala 26:23]
  wire  mem_io_em_bus_MemWen; // @[TopMain.scala 26:23]
  wire [63:0] mem_io_em_bus_Memwdata; // @[TopMain.scala 26:23]
  wire [7:0] mem_io_em_bus_wmask; // @[TopMain.scala 26:23]
  wire  mem_io_mw_bus_gr_we; // @[TopMain.scala 26:23]
  wire [4:0] mem_io_mw_bus_dest; // @[TopMain.scala 26:23]
  wire [63:0] mem_io_mw_bus_final_result; // @[TopMain.scala 26:23]
  wire [31:0] mem_io_mw_bus_mem_pc; // @[TopMain.scala 26:23]
  wire [31:0] mem_io_mw_bus_inst; // @[TopMain.scala 26:23]
  wire [63:0] mem_io_mw_bus_csr_wdata; // @[TopMain.scala 26:23]
  wire  mem_io_mw_bus_csr_wen; // @[TopMain.scala 26:23]
  wire [2:0] mem_io_mw_bus_csr_waddr1; // @[TopMain.scala 26:23]
  wire [2:0] mem_io_mw_bus_csr_waddr2; // @[TopMain.scala 26:23]
  wire  mem_io_mw_bus_eval; // @[TopMain.scala 26:23]
  wire  mem_io_ms_dest_valid_gr_we; // @[TopMain.scala 26:23]
  wire  mem_io_ms_dest_valid_ms_valid; // @[TopMain.scala 26:23]
  wire [4:0] mem_io_ms_dest_valid_dest; // @[TopMain.scala 26:23]
  wire [63:0] mem_io_ms_dest_valid_ms_forward_data; // @[TopMain.scala 26:23]
  wire  mem_io_ms_dest_valid_ms_is_ld; // @[TopMain.scala 26:23]
  wire  mem_io_ms_dest_valid_ms_to_ws_valid; // @[TopMain.scala 26:23]
  wire  mem_io_ms_dest_valid_ms_ready_go; // @[TopMain.scala 26:23]
  wire [63:0] mem_io_data_sram_rdata; // @[TopMain.scala 26:23]
  wire [63:0] mem_io_mem_result; // @[TopMain.scala 26:23]
  wire [2:0] mem_io_ld_type; // @[TopMain.scala 26:23]
  wire  mem_io_data_sram_data_ok; // @[TopMain.scala 26:23]
  wire  mem_io_data_sram_req; // @[TopMain.scala 26:23]
  wire  mem_io_data_sram_we; // @[TopMain.scala 26:23]
  wire [31:0] mem_io_data_sram_addr; // @[TopMain.scala 26:23]
  wire [63:0] mem_io_data_sram_wdata; // @[TopMain.scala 26:23]
  wire [7:0] mem_io_data_sram_wmask; // @[TopMain.scala 26:23]
  wire  mem_io_data_sram_addr_ok; // @[TopMain.scala 26:23]
  wire  wbu_clock; // @[TopMain.scala 27:23]
  wire  wbu_reset; // @[TopMain.scala 27:23]
  wire  wbu_io_ws_allowin; // @[TopMain.scala 27:23]
  wire  wbu_io_ms_to_ws_valid; // @[TopMain.scala 27:23]
  wire  wbu_io_mw_bus_gr_we; // @[TopMain.scala 27:23]
  wire [4:0] wbu_io_mw_bus_dest; // @[TopMain.scala 27:23]
  wire [63:0] wbu_io_mw_bus_final_result; // @[TopMain.scala 27:23]
  wire [31:0] wbu_io_mw_bus_mem_pc; // @[TopMain.scala 27:23]
  wire [31:0] wbu_io_mw_bus_inst; // @[TopMain.scala 27:23]
  wire [63:0] wbu_io_mw_bus_csr_wdata; // @[TopMain.scala 27:23]
  wire  wbu_io_mw_bus_csr_wen; // @[TopMain.scala 27:23]
  wire [2:0] wbu_io_mw_bus_csr_waddr1; // @[TopMain.scala 27:23]
  wire [2:0] wbu_io_mw_bus_csr_waddr2; // @[TopMain.scala 27:23]
  wire  wbu_io_mw_bus_eval; // @[TopMain.scala 27:23]
  wire  wbu_io_rf_bus_rf_we; // @[TopMain.scala 27:23]
  wire [4:0] wbu_io_rf_bus_rf_waddr; // @[TopMain.scala 27:23]
  wire [63:0] wbu_io_rf_bus_rf_wdata; // @[TopMain.scala 27:23]
  wire [31:0] wbu_io_rf_bus_wb_pc; // @[TopMain.scala 27:23]
  wire [31:0] wbu_io_rf_bus_wb_inst; // @[TopMain.scala 27:23]
  wire [63:0] wbu_io_rf_bus_csr_wdata; // @[TopMain.scala 27:23]
  wire  wbu_io_rf_bus_csr_wen; // @[TopMain.scala 27:23]
  wire [2:0] wbu_io_rf_bus_csr_waddr1; // @[TopMain.scala 27:23]
  wire [2:0] wbu_io_rf_bus_csr_waddr2; // @[TopMain.scala 27:23]
  wire  wbu_io_rf_bus_eval; // @[TopMain.scala 27:23]
  wire  wbu_io_in_WB; // @[TopMain.scala 27:23]
  wire  wbu_io_ws_dest_valid_gr_we; // @[TopMain.scala 27:23]
  wire  wbu_io_ws_dest_valid_ws_valid; // @[TopMain.scala 27:23]
  wire [4:0] wbu_io_ws_dest_valid_dest; // @[TopMain.scala 27:23]
  wire [63:0] wbu_io_ws_dest_valid_ws_forward_data; // @[TopMain.scala 27:23]
  wire [63:0] wbu_io_wb_pc; // @[TopMain.scala 27:23]
  wire [63:0] wbu_io_wb_inst; // @[TopMain.scala 27:23]
  wire [63:0] dpi_rf_0; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_1; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_2; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_3; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_4; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_5; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_6; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_7; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_8; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_9; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_10; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_11; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_12; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_13; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_14; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_15; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_16; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_17; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_18; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_19; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_20; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_21; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_22; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_23; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_24; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_25; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_26; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_27; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_28; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_29; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_30; // @[TopMain.scala 28:23]
  wire [63:0] dpi_rf_31; // @[TopMain.scala 28:23]
  wire [63:0] dpi_csr_0; // @[TopMain.scala 28:23]
  wire [63:0] dpi_csr_1; // @[TopMain.scala 28:23]
  wire [63:0] dpi_csr_2; // @[TopMain.scala 28:23]
  wire [63:0] dpi_csr_3; // @[TopMain.scala 28:23]
  wire [63:0] dpi_csr_4; // @[TopMain.scala 28:23]
  wire [31:0] dpi_inst; // @[TopMain.scala 28:23]
  wire [63:0] dpi_pc; // @[TopMain.scala 28:23]
  wire [31:0] dpi_eval; // @[TopMain.scala 28:23]
  wire  axi_clock; // @[TopMain.scala 29:23]
  wire  axi_reset; // @[TopMain.scala 29:23]
  wire [3:0] axi_io_arid; // @[TopMain.scala 29:23]
  wire [63:0] axi_io_araddr; // @[TopMain.scala 29:23]
  wire  axi_io_arvalid; // @[TopMain.scala 29:23]
  wire  axi_io_arready; // @[TopMain.scala 29:23]
  wire [63:0] axi_io_rdata; // @[TopMain.scala 29:23]
  wire [127:0] axi_io_icache_rdata; // @[TopMain.scala 29:23]
  wire  axi_io_rvalid; // @[TopMain.scala 29:23]
  wire  axi_io_rready; // @[TopMain.scala 29:23]
  wire [63:0] axi_io_awaddr; // @[TopMain.scala 29:23]
  wire  axi_io_awvalid; // @[TopMain.scala 29:23]
  wire  axi_io_awready; // @[TopMain.scala 29:23]
  wire [63:0] axi_io_wdata; // @[TopMain.scala 29:23]
  wire [7:0] axi_io_wstrb; // @[TopMain.scala 29:23]
  wire  axi_io_wvalid; // @[TopMain.scala 29:23]
  wire  axi_io_wready; // @[TopMain.scala 29:23]
  wire  axi_io_bvalid; // @[TopMain.scala 29:23]
  wire  axi_io_bready; // @[TopMain.scala 29:23]
  wire  axi_io_inst_sram_req; // @[TopMain.scala 29:23]
  wire [63:0] axi_io_inst_sram_addr; // @[TopMain.scala 29:23]
  wire [127:0] axi_io_inst_sram_rdata; // @[TopMain.scala 29:23]
  wire  axi_io_inst_sram_addr_ok; // @[TopMain.scala 29:23]
  wire  axi_io_inst_sram_data_ok; // @[TopMain.scala 29:23]
  wire  axi_io_data_sram_req; // @[TopMain.scala 29:23]
  wire  axi_io_data_sram_wr; // @[TopMain.scala 29:23]
  wire [7:0] axi_io_data_sram_wstrb; // @[TopMain.scala 29:23]
  wire [63:0] axi_io_data_sram_addr; // @[TopMain.scala 29:23]
  wire [63:0] axi_io_data_sram_wdata; // @[TopMain.scala 29:23]
  wire [63:0] axi_io_data_sram_rdata; // @[TopMain.scala 29:23]
  wire  axi_io_data_sram_addr_ok; // @[TopMain.scala 29:23]
  wire  axi_io_data_sram_data_ok; // @[TopMain.scala 29:23]
  wire  axi_mem_reset; // @[TopMain.scala 30:23]
  wire  axi_mem_clock; // @[TopMain.scala 30:23]
  wire [3:0] axi_mem_arid; // @[TopMain.scala 30:23]
  wire [63:0] axi_mem_araddr; // @[TopMain.scala 30:23]
  wire  axi_mem_arvalid; // @[TopMain.scala 30:23]
  wire  axi_mem_arready; // @[TopMain.scala 30:23]
  wire [63:0] axi_mem_rdata; // @[TopMain.scala 30:23]
  wire [127:0] axi_mem_icache_rdata; // @[TopMain.scala 30:23]
  wire  axi_mem_rvalid; // @[TopMain.scala 30:23]
  wire  axi_mem_rready; // @[TopMain.scala 30:23]
  wire [3:0] axi_mem_awid; // @[TopMain.scala 30:23]
  wire [63:0] axi_mem_awaddr; // @[TopMain.scala 30:23]
  wire  axi_mem_awvalid; // @[TopMain.scala 30:23]
  wire  axi_mem_awready; // @[TopMain.scala 30:23]
  wire [63:0] axi_mem_wdata; // @[TopMain.scala 30:23]
  wire [7:0] axi_mem_wstrb; // @[TopMain.scala 30:23]
  wire  axi_mem_wvalid; // @[TopMain.scala 30:23]
  wire  axi_mem_wready; // @[TopMain.scala 30:23]
  wire  axi_mem_bvalid; // @[TopMain.scala 30:23]
  wire  axi_mem_bready; // @[TopMain.scala 30:23]
  wire  icache_clock; // @[TopMain.scala 31:24]
  wire  icache_reset; // @[TopMain.scala 31:24]
  wire  icache_io_valid; // @[TopMain.scala 31:24]
  wire [63:0] icache_io_addr; // @[TopMain.scala 31:24]
  wire [63:0] icache_io_rdata; // @[TopMain.scala 31:24]
  wire  icache_io_addr_ok; // @[TopMain.scala 31:24]
  wire  icache_io_data_ok; // @[TopMain.scala 31:24]
  wire  icache_io_rd_req; // @[TopMain.scala 31:24]
  wire [31:0] icache_io_rd_addr; // @[TopMain.scala 31:24]
  wire  icache_io_rd_rdy; // @[TopMain.scala 31:24]
  wire [127:0] icache_io_rd_data; // @[TopMain.scala 31:24]
  wire  icache_io_inst_sram_data_ok; // @[TopMain.scala 31:24]
  IFU ifu ( // @[TopMain.scala 23:23]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_reset(ifu_io_reset),
    .io_fd_bus_inst(ifu_io_fd_bus_inst),
    .io_fd_bus_pc(ifu_io_fd_bus_pc),
    .io_ds_allowin(ifu_io_ds_allowin),
    .io_fs_to_ds_valid(ifu_io_fs_to_ds_valid),
    .io_br_bus_br_taken(ifu_io_br_bus_br_taken),
    .io_br_bus_br_target(ifu_io_br_bus_br_target),
    .io_br_bus_rawblock(ifu_io_br_bus_rawblock),
    .io_br_bus_csr_rdata(ifu_io_br_bus_csr_rdata),
    .io_br_bus_eval(ifu_io_br_bus_eval),
    .io_br_bus_mret(ifu_io_br_bus_mret),
    .io_inst_sram_req(ifu_io_inst_sram_req),
    .io_inst_sram_addr(ifu_io_inst_sram_addr),
    .io_inst_sram_rdata(ifu_io_inst_sram_rdata),
    .io_inst_sram_addr_ok(ifu_io_inst_sram_addr_ok),
    .io_inst_sram_data_ok(ifu_io_inst_sram_data_ok)
  );
  IDU idu ( // @[TopMain.scala 24:23]
    .clock(idu_clock),
    .reset(idu_reset),
    .io_es_allowin(idu_io_es_allowin),
    .io_ds_allowin(idu_io_ds_allowin),
    .io_fs_to_ds_valid(idu_io_fs_to_ds_valid),
    .io_ds_to_es_valid(idu_io_ds_to_es_valid),
    .io_fd_bus_inst(idu_io_fd_bus_inst),
    .io_fd_bus_pc(idu_io_fd_bus_pc),
    .io_de_bus_OP(idu_io_de_bus_OP),
    .io_de_bus_res_from_mem(idu_io_de_bus_res_from_mem),
    .io_de_bus_gr_we(idu_io_de_bus_gr_we),
    .io_de_bus_MemWen(idu_io_de_bus_MemWen),
    .io_de_bus_wmask(idu_io_de_bus_wmask),
    .io_de_bus_ds_pc(idu_io_de_bus_ds_pc),
    .io_de_bus_dest(idu_io_de_bus_dest),
    .io_de_bus_imm(idu_io_de_bus_imm),
    .io_de_bus_rdata1(idu_io_de_bus_rdata1),
    .io_de_bus_rdata2(idu_io_de_bus_rdata2),
    .io_de_bus_ld_type(idu_io_de_bus_ld_type),
    .io_de_bus_inst(idu_io_de_bus_inst),
    .io_de_bus_csr_rdata(idu_io_de_bus_csr_rdata),
    .io_de_bus_csr_waddr1(idu_io_de_bus_csr_waddr1),
    .io_de_bus_csr_waddr2(idu_io_de_bus_csr_waddr2),
    .io_de_bus_csr_raddr(idu_io_de_bus_csr_raddr),
    .io_de_bus_csr_ren(idu_io_de_bus_csr_ren),
    .io_de_bus_csr_wen(idu_io_de_bus_csr_wen),
    .io_de_bus_eval(idu_io_de_bus_eval),
    .io_de_bus_is_ld(idu_io_de_bus_is_ld),
    .io_br_bus_br_taken(idu_io_br_bus_br_taken),
    .io_br_bus_br_target(idu_io_br_bus_br_target),
    .io_br_bus_rawblock(idu_io_br_bus_rawblock),
    .io_br_bus_csr_rdata(idu_io_br_bus_csr_rdata),
    .io_br_bus_eval(idu_io_br_bus_eval),
    .io_br_bus_mret(idu_io_br_bus_mret),
    .io_rf_bus_rf_we(idu_io_rf_bus_rf_we),
    .io_rf_bus_rf_waddr(idu_io_rf_bus_rf_waddr),
    .io_rf_bus_rf_wdata(idu_io_rf_bus_rf_wdata),
    .io_rf_bus_wb_pc(idu_io_rf_bus_wb_pc),
    .io_rf_bus_wb_inst(idu_io_rf_bus_wb_inst),
    .io_rf_bus_csr_wdata(idu_io_rf_bus_csr_wdata),
    .io_rf_bus_csr_wen(idu_io_rf_bus_csr_wen),
    .io_rf_bus_csr_waddr1(idu_io_rf_bus_csr_waddr1),
    .io_rf_bus_csr_waddr2(idu_io_rf_bus_csr_waddr2),
    .io_rf_bus_eval(idu_io_rf_bus_eval),
    .io_es_dest_valid_gr_we(idu_io_es_dest_valid_gr_we),
    .io_es_dest_valid_es_valid(idu_io_es_dest_valid_es_valid),
    .io_es_dest_valid_dest(idu_io_es_dest_valid_dest),
    .io_es_dest_valid_es_forward_data(idu_io_es_dest_valid_es_forward_data),
    .io_es_dest_valid_es_is_ld(idu_io_es_dest_valid_es_is_ld),
    .io_es_dest_valid_es_ready_go(idu_io_es_dest_valid_es_ready_go),
    .io_es_dest_valid_es_to_ms_valid(idu_io_es_dest_valid_es_to_ms_valid),
    .io_ms_dest_valid_gr_we(idu_io_ms_dest_valid_gr_we),
    .io_ms_dest_valid_ms_valid(idu_io_ms_dest_valid_ms_valid),
    .io_ms_dest_valid_dest(idu_io_ms_dest_valid_dest),
    .io_ms_dest_valid_ms_forward_data(idu_io_ms_dest_valid_ms_forward_data),
    .io_ms_dest_valid_ms_is_ld(idu_io_ms_dest_valid_ms_is_ld),
    .io_ms_dest_valid_ms_to_ws_valid(idu_io_ms_dest_valid_ms_to_ws_valid),
    .io_ms_dest_valid_ms_ready_go(idu_io_ms_dest_valid_ms_ready_go),
    .io_ws_dest_valid_gr_we(idu_io_ws_dest_valid_gr_we),
    .io_ws_dest_valid_ws_valid(idu_io_ws_dest_valid_ws_valid),
    .io_ws_dest_valid_dest(idu_io_ws_dest_valid_dest),
    .io_ws_dest_valid_ws_forward_data(idu_io_ws_dest_valid_ws_forward_data)
  );
  EXU exu ( // @[TopMain.scala 25:23]
    .clock(exu_clock),
    .reset(exu_reset),
    .io_ms_allowin(exu_io_ms_allowin),
    .io_es_allowin(exu_io_es_allowin),
    .io_ds_to_es_valid(exu_io_ds_to_es_valid),
    .io_es_to_ms_valid(exu_io_es_to_ms_valid),
    .io_de_bus_OP(exu_io_de_bus_OP),
    .io_de_bus_res_from_mem(exu_io_de_bus_res_from_mem),
    .io_de_bus_gr_we(exu_io_de_bus_gr_we),
    .io_de_bus_MemWen(exu_io_de_bus_MemWen),
    .io_de_bus_wmask(exu_io_de_bus_wmask),
    .io_de_bus_ds_pc(exu_io_de_bus_ds_pc),
    .io_de_bus_dest(exu_io_de_bus_dest),
    .io_de_bus_imm(exu_io_de_bus_imm),
    .io_de_bus_rdata1(exu_io_de_bus_rdata1),
    .io_de_bus_rdata2(exu_io_de_bus_rdata2),
    .io_de_bus_ld_type(exu_io_de_bus_ld_type),
    .io_de_bus_inst(exu_io_de_bus_inst),
    .io_de_bus_csr_rdata(exu_io_de_bus_csr_rdata),
    .io_de_bus_csr_waddr1(exu_io_de_bus_csr_waddr1),
    .io_de_bus_csr_waddr2(exu_io_de_bus_csr_waddr2),
    .io_de_bus_csr_wen(exu_io_de_bus_csr_wen),
    .io_de_bus_eval(exu_io_de_bus_eval),
    .io_de_bus_is_ld(exu_io_de_bus_is_ld),
    .io_em_bus_res_from_mem(exu_io_em_bus_res_from_mem),
    .io_em_bus_gr_we(exu_io_em_bus_gr_we),
    .io_em_bus_dest(exu_io_em_bus_dest),
    .io_em_bus_alu_result(exu_io_em_bus_alu_result),
    .io_em_bus_ex_pc(exu_io_em_bus_ex_pc),
    .io_em_bus_ld_type(exu_io_em_bus_ld_type),
    .io_em_bus_inst(exu_io_em_bus_inst),
    .io_em_bus_csr_wdata(exu_io_em_bus_csr_wdata),
    .io_em_bus_csr_wen(exu_io_em_bus_csr_wen),
    .io_em_bus_csr_waddr1(exu_io_em_bus_csr_waddr1),
    .io_em_bus_csr_waddr2(exu_io_em_bus_csr_waddr2),
    .io_em_bus_eval(exu_io_em_bus_eval),
    .io_em_bus_is_ld(exu_io_em_bus_is_ld),
    .io_em_bus_MemWen(exu_io_em_bus_MemWen),
    .io_em_bus_Memwdata(exu_io_em_bus_Memwdata),
    .io_em_bus_wmask(exu_io_em_bus_wmask),
    .io_es_dest_valid_gr_we(exu_io_es_dest_valid_gr_we),
    .io_es_dest_valid_es_valid(exu_io_es_dest_valid_es_valid),
    .io_es_dest_valid_dest(exu_io_es_dest_valid_dest),
    .io_es_dest_valid_es_forward_data(exu_io_es_dest_valid_es_forward_data),
    .io_es_dest_valid_es_is_ld(exu_io_es_dest_valid_es_is_ld),
    .io_es_dest_valid_es_ready_go(exu_io_es_dest_valid_es_ready_go),
    .io_es_dest_valid_es_to_ms_valid(exu_io_es_dest_valid_es_to_ms_valid)
  );
  MEM mem ( // @[TopMain.scala 26:23]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_ms_allowin(mem_io_ms_allowin),
    .io_es_to_ms_valid(mem_io_es_to_ms_valid),
    .io_ms_to_ws_valid(mem_io_ms_to_ws_valid),
    .io_em_bus_res_from_mem(mem_io_em_bus_res_from_mem),
    .io_em_bus_gr_we(mem_io_em_bus_gr_we),
    .io_em_bus_dest(mem_io_em_bus_dest),
    .io_em_bus_alu_result(mem_io_em_bus_alu_result),
    .io_em_bus_ex_pc(mem_io_em_bus_ex_pc),
    .io_em_bus_ld_type(mem_io_em_bus_ld_type),
    .io_em_bus_inst(mem_io_em_bus_inst),
    .io_em_bus_csr_wdata(mem_io_em_bus_csr_wdata),
    .io_em_bus_csr_wen(mem_io_em_bus_csr_wen),
    .io_em_bus_csr_waddr1(mem_io_em_bus_csr_waddr1),
    .io_em_bus_csr_waddr2(mem_io_em_bus_csr_waddr2),
    .io_em_bus_eval(mem_io_em_bus_eval),
    .io_em_bus_is_ld(mem_io_em_bus_is_ld),
    .io_em_bus_MemWen(mem_io_em_bus_MemWen),
    .io_em_bus_Memwdata(mem_io_em_bus_Memwdata),
    .io_em_bus_wmask(mem_io_em_bus_wmask),
    .io_mw_bus_gr_we(mem_io_mw_bus_gr_we),
    .io_mw_bus_dest(mem_io_mw_bus_dest),
    .io_mw_bus_final_result(mem_io_mw_bus_final_result),
    .io_mw_bus_mem_pc(mem_io_mw_bus_mem_pc),
    .io_mw_bus_inst(mem_io_mw_bus_inst),
    .io_mw_bus_csr_wdata(mem_io_mw_bus_csr_wdata),
    .io_mw_bus_csr_wen(mem_io_mw_bus_csr_wen),
    .io_mw_bus_csr_waddr1(mem_io_mw_bus_csr_waddr1),
    .io_mw_bus_csr_waddr2(mem_io_mw_bus_csr_waddr2),
    .io_mw_bus_eval(mem_io_mw_bus_eval),
    .io_ms_dest_valid_gr_we(mem_io_ms_dest_valid_gr_we),
    .io_ms_dest_valid_ms_valid(mem_io_ms_dest_valid_ms_valid),
    .io_ms_dest_valid_dest(mem_io_ms_dest_valid_dest),
    .io_ms_dest_valid_ms_forward_data(mem_io_ms_dest_valid_ms_forward_data),
    .io_ms_dest_valid_ms_is_ld(mem_io_ms_dest_valid_ms_is_ld),
    .io_ms_dest_valid_ms_to_ws_valid(mem_io_ms_dest_valid_ms_to_ws_valid),
    .io_ms_dest_valid_ms_ready_go(mem_io_ms_dest_valid_ms_ready_go),
    .io_data_sram_rdata(mem_io_data_sram_rdata),
    .io_mem_result(mem_io_mem_result),
    .io_ld_type(mem_io_ld_type),
    .io_data_sram_data_ok(mem_io_data_sram_data_ok),
    .io_data_sram_req(mem_io_data_sram_req),
    .io_data_sram_we(mem_io_data_sram_we),
    .io_data_sram_addr(mem_io_data_sram_addr),
    .io_data_sram_wdata(mem_io_data_sram_wdata),
    .io_data_sram_wmask(mem_io_data_sram_wmask),
    .io_data_sram_addr_ok(mem_io_data_sram_addr_ok)
  );
  WBU wbu ( // @[TopMain.scala 27:23]
    .clock(wbu_clock),
    .reset(wbu_reset),
    .io_ws_allowin(wbu_io_ws_allowin),
    .io_ms_to_ws_valid(wbu_io_ms_to_ws_valid),
    .io_mw_bus_gr_we(wbu_io_mw_bus_gr_we),
    .io_mw_bus_dest(wbu_io_mw_bus_dest),
    .io_mw_bus_final_result(wbu_io_mw_bus_final_result),
    .io_mw_bus_mem_pc(wbu_io_mw_bus_mem_pc),
    .io_mw_bus_inst(wbu_io_mw_bus_inst),
    .io_mw_bus_csr_wdata(wbu_io_mw_bus_csr_wdata),
    .io_mw_bus_csr_wen(wbu_io_mw_bus_csr_wen),
    .io_mw_bus_csr_waddr1(wbu_io_mw_bus_csr_waddr1),
    .io_mw_bus_csr_waddr2(wbu_io_mw_bus_csr_waddr2),
    .io_mw_bus_eval(wbu_io_mw_bus_eval),
    .io_rf_bus_rf_we(wbu_io_rf_bus_rf_we),
    .io_rf_bus_rf_waddr(wbu_io_rf_bus_rf_waddr),
    .io_rf_bus_rf_wdata(wbu_io_rf_bus_rf_wdata),
    .io_rf_bus_wb_pc(wbu_io_rf_bus_wb_pc),
    .io_rf_bus_wb_inst(wbu_io_rf_bus_wb_inst),
    .io_rf_bus_csr_wdata(wbu_io_rf_bus_csr_wdata),
    .io_rf_bus_csr_wen(wbu_io_rf_bus_csr_wen),
    .io_rf_bus_csr_waddr1(wbu_io_rf_bus_csr_waddr1),
    .io_rf_bus_csr_waddr2(wbu_io_rf_bus_csr_waddr2),
    .io_rf_bus_eval(wbu_io_rf_bus_eval),
    .io_in_WB(wbu_io_in_WB),
    .io_ws_dest_valid_gr_we(wbu_io_ws_dest_valid_gr_we),
    .io_ws_dest_valid_ws_valid(wbu_io_ws_dest_valid_ws_valid),
    .io_ws_dest_valid_dest(wbu_io_ws_dest_valid_dest),
    .io_ws_dest_valid_ws_forward_data(wbu_io_ws_dest_valid_ws_forward_data),
    .io_wb_pc(wbu_io_wb_pc),
    .io_wb_inst(wbu_io_wb_inst)
  );
  DPI dpi ( // @[TopMain.scala 28:23]
    .rf_0(dpi_rf_0),
    .rf_1(dpi_rf_1),
    .rf_2(dpi_rf_2),
    .rf_3(dpi_rf_3),
    .rf_4(dpi_rf_4),
    .rf_5(dpi_rf_5),
    .rf_6(dpi_rf_6),
    .rf_7(dpi_rf_7),
    .rf_8(dpi_rf_8),
    .rf_9(dpi_rf_9),
    .rf_10(dpi_rf_10),
    .rf_11(dpi_rf_11),
    .rf_12(dpi_rf_12),
    .rf_13(dpi_rf_13),
    .rf_14(dpi_rf_14),
    .rf_15(dpi_rf_15),
    .rf_16(dpi_rf_16),
    .rf_17(dpi_rf_17),
    .rf_18(dpi_rf_18),
    .rf_19(dpi_rf_19),
    .rf_20(dpi_rf_20),
    .rf_21(dpi_rf_21),
    .rf_22(dpi_rf_22),
    .rf_23(dpi_rf_23),
    .rf_24(dpi_rf_24),
    .rf_25(dpi_rf_25),
    .rf_26(dpi_rf_26),
    .rf_27(dpi_rf_27),
    .rf_28(dpi_rf_28),
    .rf_29(dpi_rf_29),
    .rf_30(dpi_rf_30),
    .rf_31(dpi_rf_31),
    .csr_0(dpi_csr_0),
    .csr_1(dpi_csr_1),
    .csr_2(dpi_csr_2),
    .csr_3(dpi_csr_3),
    .csr_4(dpi_csr_4),
    .inst(dpi_inst),
    .pc(dpi_pc),
    .eval(dpi_eval)
  );
  AXI axi ( // @[TopMain.scala 29:23]
    .clock(axi_clock),
    .reset(axi_reset),
    .io_arid(axi_io_arid),
    .io_araddr(axi_io_araddr),
    .io_arvalid(axi_io_arvalid),
    .io_arready(axi_io_arready),
    .io_rdata(axi_io_rdata),
    .io_icache_rdata(axi_io_icache_rdata),
    .io_rvalid(axi_io_rvalid),
    .io_rready(axi_io_rready),
    .io_awaddr(axi_io_awaddr),
    .io_awvalid(axi_io_awvalid),
    .io_awready(axi_io_awready),
    .io_wdata(axi_io_wdata),
    .io_wstrb(axi_io_wstrb),
    .io_wvalid(axi_io_wvalid),
    .io_wready(axi_io_wready),
    .io_bvalid(axi_io_bvalid),
    .io_bready(axi_io_bready),
    .io_inst_sram_req(axi_io_inst_sram_req),
    .io_inst_sram_addr(axi_io_inst_sram_addr),
    .io_inst_sram_rdata(axi_io_inst_sram_rdata),
    .io_inst_sram_addr_ok(axi_io_inst_sram_addr_ok),
    .io_inst_sram_data_ok(axi_io_inst_sram_data_ok),
    .io_data_sram_req(axi_io_data_sram_req),
    .io_data_sram_wr(axi_io_data_sram_wr),
    .io_data_sram_wstrb(axi_io_data_sram_wstrb),
    .io_data_sram_addr(axi_io_data_sram_addr),
    .io_data_sram_wdata(axi_io_data_sram_wdata),
    .io_data_sram_rdata(axi_io_data_sram_rdata),
    .io_data_sram_addr_ok(axi_io_data_sram_addr_ok),
    .io_data_sram_data_ok(axi_io_data_sram_data_ok)
  );
  AXI_mem axi_mem ( // @[TopMain.scala 30:23]
    .reset(axi_mem_reset),
    .clock(axi_mem_clock),
    .arid(axi_mem_arid),
    .araddr(axi_mem_araddr),
    .arvalid(axi_mem_arvalid),
    .arready(axi_mem_arready),
    .rdata(axi_mem_rdata),
    .icache_rdata(axi_mem_icache_rdata),
    .rvalid(axi_mem_rvalid),
    .rready(axi_mem_rready),
    .awid(axi_mem_awid),
    .awaddr(axi_mem_awaddr),
    .awvalid(axi_mem_awvalid),
    .awready(axi_mem_awready),
    .wdata(axi_mem_wdata),
    .wstrb(axi_mem_wstrb),
    .wvalid(axi_mem_wvalid),
    .wready(axi_mem_wready),
    .bvalid(axi_mem_bvalid),
    .bready(axi_mem_bready)
  );
  icache icache ( // @[TopMain.scala 31:24]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_valid(icache_io_valid),
    .io_addr(icache_io_addr),
    .io_rdata(icache_io_rdata),
    .io_addr_ok(icache_io_addr_ok),
    .io_data_ok(icache_io_data_ok),
    .io_rd_req(icache_io_rd_req),
    .io_rd_addr(icache_io_rd_addr),
    .io_rd_rdy(icache_io_rd_rdy),
    .io_rd_data(icache_io_rd_data),
    .io_inst_sram_data_ok(icache_io_inst_sram_data_ok)
  );
  assign io_fs_pc = ifu_io_fd_bus_pc; // @[TopMain.scala 85:17]
  assign io_op = idu_io_de_bus_OP[6:0]; // @[TopMain.scala 86:17]
  assign io_in_WB = wbu_io_in_WB; // @[TopMain.scala 87:17]
  assign io_wb_pc = wbu_io_wb_pc[31:0]; // @[TopMain.scala 88:17]
  assign io_wb_inst = wbu_io_wb_inst[31:0]; // @[TopMain.scala 89:17]
  assign io_ds_pc = idu_io_de_bus_ds_pc; // @[TopMain.scala 90:17]
  assign io_mem_result = mem_io_mem_result; // @[TopMain.scala 91:17]
  assign io_ld_type = mem_io_ld_type; // @[TopMain.scala 92:17]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_reset = reset; // @[TopMain.scala 35:16]
  assign ifu_io_ds_allowin = idu_io_ds_allowin; // @[TopMain.scala 36:21]
  assign ifu_io_br_bus_br_taken = idu_io_br_bus_br_taken; // @[TopMain.scala 37:17]
  assign ifu_io_br_bus_br_target = idu_io_br_bus_br_target; // @[TopMain.scala 37:17]
  assign ifu_io_br_bus_rawblock = idu_io_br_bus_rawblock; // @[TopMain.scala 37:17]
  assign ifu_io_br_bus_csr_rdata = idu_io_br_bus_csr_rdata; // @[TopMain.scala 37:17]
  assign ifu_io_br_bus_eval = idu_io_br_bus_eval; // @[TopMain.scala 37:17]
  assign ifu_io_br_bus_mret = idu_io_br_bus_mret; // @[TopMain.scala 37:17]
  assign ifu_io_inst_sram_rdata = icache_io_rdata; // @[TopMain.scala 38:26]
  assign ifu_io_inst_sram_addr_ok = icache_io_addr_ok; // @[TopMain.scala 40:28]
  assign ifu_io_inst_sram_data_ok = icache_io_data_ok; // @[TopMain.scala 39:28]
  assign idu_clock = clock;
  assign idu_reset = reset;
  assign idu_io_es_allowin = exu_io_es_allowin; // @[TopMain.scala 51:21]
  assign idu_io_fs_to_ds_valid = ifu_io_fs_to_ds_valid; // @[TopMain.scala 52:25]
  assign idu_io_fd_bus_inst = ifu_io_fd_bus_inst; // @[TopMain.scala 53:17]
  assign idu_io_fd_bus_pc = ifu_io_fd_bus_pc; // @[TopMain.scala 53:17]
  assign idu_io_rf_bus_rf_we = wbu_io_rf_bus_rf_we; // @[TopMain.scala 54:17]
  assign idu_io_rf_bus_rf_waddr = wbu_io_rf_bus_rf_waddr; // @[TopMain.scala 54:17]
  assign idu_io_rf_bus_rf_wdata = wbu_io_rf_bus_rf_wdata; // @[TopMain.scala 54:17]
  assign idu_io_rf_bus_wb_pc = wbu_io_rf_bus_wb_pc; // @[TopMain.scala 54:17]
  assign idu_io_rf_bus_wb_inst = wbu_io_rf_bus_wb_inst; // @[TopMain.scala 54:17]
  assign idu_io_rf_bus_csr_wdata = wbu_io_rf_bus_csr_wdata; // @[TopMain.scala 54:17]
  assign idu_io_rf_bus_csr_wen = wbu_io_rf_bus_csr_wen; // @[TopMain.scala 54:17]
  assign idu_io_rf_bus_csr_waddr1 = wbu_io_rf_bus_csr_waddr1; // @[TopMain.scala 54:17]
  assign idu_io_rf_bus_csr_waddr2 = wbu_io_rf_bus_csr_waddr2; // @[TopMain.scala 54:17]
  assign idu_io_rf_bus_eval = wbu_io_rf_bus_eval; // @[TopMain.scala 54:17]
  assign idu_io_es_dest_valid_gr_we = exu_io_es_dest_valid_gr_we; // @[TopMain.scala 55:24]
  assign idu_io_es_dest_valid_es_valid = exu_io_es_dest_valid_es_valid; // @[TopMain.scala 55:24]
  assign idu_io_es_dest_valid_dest = exu_io_es_dest_valid_dest; // @[TopMain.scala 55:24]
  assign idu_io_es_dest_valid_es_forward_data = exu_io_es_dest_valid_es_forward_data; // @[TopMain.scala 55:24]
  assign idu_io_es_dest_valid_es_is_ld = exu_io_es_dest_valid_es_is_ld; // @[TopMain.scala 55:24]
  assign idu_io_es_dest_valid_es_ready_go = exu_io_es_dest_valid_es_ready_go; // @[TopMain.scala 55:24]
  assign idu_io_es_dest_valid_es_to_ms_valid = exu_io_es_dest_valid_es_to_ms_valid; // @[TopMain.scala 55:24]
  assign idu_io_ms_dest_valid_gr_we = mem_io_ms_dest_valid_gr_we; // @[TopMain.scala 56:24]
  assign idu_io_ms_dest_valid_ms_valid = mem_io_ms_dest_valid_ms_valid; // @[TopMain.scala 56:24]
  assign idu_io_ms_dest_valid_dest = mem_io_ms_dest_valid_dest; // @[TopMain.scala 56:24]
  assign idu_io_ms_dest_valid_ms_forward_data = mem_io_ms_dest_valid_ms_forward_data; // @[TopMain.scala 56:24]
  assign idu_io_ms_dest_valid_ms_is_ld = mem_io_ms_dest_valid_ms_is_ld; // @[TopMain.scala 56:24]
  assign idu_io_ms_dest_valid_ms_to_ws_valid = mem_io_ms_dest_valid_ms_to_ws_valid; // @[TopMain.scala 56:24]
  assign idu_io_ms_dest_valid_ms_ready_go = mem_io_ms_dest_valid_ms_ready_go; // @[TopMain.scala 56:24]
  assign idu_io_ws_dest_valid_gr_we = wbu_io_ws_dest_valid_gr_we; // @[TopMain.scala 57:24]
  assign idu_io_ws_dest_valid_ws_valid = wbu_io_ws_dest_valid_ws_valid; // @[TopMain.scala 57:24]
  assign idu_io_ws_dest_valid_dest = wbu_io_ws_dest_valid_dest; // @[TopMain.scala 57:24]
  assign idu_io_ws_dest_valid_ws_forward_data = wbu_io_ws_dest_valid_ws_forward_data; // @[TopMain.scala 57:24]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io_ms_allowin = mem_io_ms_allowin; // @[TopMain.scala 61:21]
  assign exu_io_ds_to_es_valid = idu_io_ds_to_es_valid; // @[TopMain.scala 62:25]
  assign exu_io_de_bus_OP = idu_io_de_bus_OP; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_res_from_mem = idu_io_de_bus_res_from_mem; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_gr_we = idu_io_de_bus_gr_we; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_MemWen = idu_io_de_bus_MemWen; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_wmask = idu_io_de_bus_wmask; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_ds_pc = idu_io_de_bus_ds_pc; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_dest = idu_io_de_bus_dest; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_imm = idu_io_de_bus_imm; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_rdata1 = idu_io_de_bus_rdata1; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_rdata2 = idu_io_de_bus_rdata2; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_ld_type = idu_io_de_bus_ld_type; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_inst = idu_io_de_bus_inst; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_csr_rdata = idu_io_de_bus_csr_rdata; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_csr_waddr1 = idu_io_de_bus_csr_waddr1; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_csr_waddr2 = idu_io_de_bus_csr_waddr2; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_csr_wen = idu_io_de_bus_csr_wen; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_eval = idu_io_de_bus_eval; // @[TopMain.scala 63:17]
  assign exu_io_de_bus_is_ld = idu_io_de_bus_is_ld; // @[TopMain.scala 63:17]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_es_to_ms_valid = exu_io_es_to_ms_valid; // @[TopMain.scala 67:25]
  assign mem_io_em_bus_res_from_mem = exu_io_em_bus_res_from_mem; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_gr_we = exu_io_em_bus_gr_we; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_dest = exu_io_em_bus_dest; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_alu_result = exu_io_em_bus_alu_result; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_ex_pc = exu_io_em_bus_ex_pc; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_ld_type = exu_io_em_bus_ld_type; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_inst = exu_io_em_bus_inst; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_csr_wdata = exu_io_em_bus_csr_wdata; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_csr_wen = exu_io_em_bus_csr_wen; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_csr_waddr1 = exu_io_em_bus_csr_waddr1; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_csr_waddr2 = exu_io_em_bus_csr_waddr2; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_eval = exu_io_em_bus_eval; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_is_ld = exu_io_em_bus_is_ld; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_MemWen = exu_io_em_bus_MemWen; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_Memwdata = exu_io_em_bus_Memwdata; // @[TopMain.scala 68:17]
  assign mem_io_em_bus_wmask = exu_io_em_bus_wmask; // @[TopMain.scala 68:17]
  assign mem_io_data_sram_rdata = axi_io_data_sram_rdata; // @[TopMain.scala 70:26]
  assign mem_io_data_sram_data_ok = axi_io_data_sram_data_ok; // @[TopMain.scala 69:28]
  assign mem_io_data_sram_addr_ok = axi_io_data_sram_addr_ok; // @[TopMain.scala 71:28]
  assign wbu_clock = clock;
  assign wbu_reset = reset;
  assign wbu_io_ms_to_ws_valid = mem_io_ms_to_ws_valid; // @[TopMain.scala 81:25]
  assign wbu_io_mw_bus_gr_we = mem_io_mw_bus_gr_we; // @[TopMain.scala 82:17]
  assign wbu_io_mw_bus_dest = mem_io_mw_bus_dest; // @[TopMain.scala 82:17]
  assign wbu_io_mw_bus_final_result = mem_io_mw_bus_final_result; // @[TopMain.scala 82:17]
  assign wbu_io_mw_bus_mem_pc = mem_io_mw_bus_mem_pc; // @[TopMain.scala 82:17]
  assign wbu_io_mw_bus_inst = mem_io_mw_bus_inst; // @[TopMain.scala 82:17]
  assign wbu_io_mw_bus_csr_wdata = mem_io_mw_bus_csr_wdata; // @[TopMain.scala 82:17]
  assign wbu_io_mw_bus_csr_wen = mem_io_mw_bus_csr_wen; // @[TopMain.scala 82:17]
  assign wbu_io_mw_bus_csr_waddr1 = mem_io_mw_bus_csr_waddr1; // @[TopMain.scala 82:17]
  assign wbu_io_mw_bus_csr_waddr2 = mem_io_mw_bus_csr_waddr2; // @[TopMain.scala 82:17]
  assign wbu_io_mw_bus_eval = mem_io_mw_bus_eval; // @[TopMain.scala 82:17]
  assign dpi_rf_0 = 64'h0;
  assign dpi_rf_1 = 64'h0;
  assign dpi_rf_2 = 64'h0;
  assign dpi_rf_3 = 64'h0;
  assign dpi_rf_4 = 64'h0;
  assign dpi_rf_5 = 64'h0;
  assign dpi_rf_6 = 64'h0;
  assign dpi_rf_7 = 64'h0;
  assign dpi_rf_8 = 64'h0;
  assign dpi_rf_9 = 64'h0;
  assign dpi_rf_10 = 64'h0;
  assign dpi_rf_11 = 64'h0;
  assign dpi_rf_12 = 64'h0;
  assign dpi_rf_13 = 64'h0;
  assign dpi_rf_14 = 64'h0;
  assign dpi_rf_15 = 64'h0;
  assign dpi_rf_16 = 64'h0;
  assign dpi_rf_17 = 64'h0;
  assign dpi_rf_18 = 64'h0;
  assign dpi_rf_19 = 64'h0;
  assign dpi_rf_20 = 64'h0;
  assign dpi_rf_21 = 64'h0;
  assign dpi_rf_22 = 64'h0;
  assign dpi_rf_23 = 64'h0;
  assign dpi_rf_24 = 64'h0;
  assign dpi_rf_25 = 64'h0;
  assign dpi_rf_26 = 64'h0;
  assign dpi_rf_27 = 64'h0;
  assign dpi_rf_28 = 64'h0;
  assign dpi_rf_29 = 64'h0;
  assign dpi_rf_30 = 64'h0;
  assign dpi_rf_31 = 64'h0;
  assign dpi_csr_0 = 64'h0;
  assign dpi_csr_1 = 64'h0;
  assign dpi_csr_2 = 64'h0;
  assign dpi_csr_3 = 64'h0;
  assign dpi_csr_4 = 64'h0;
  assign dpi_inst = 32'h0;
  assign dpi_pc = 64'h0;
  assign dpi_eval = 32'h0;
  assign axi_clock = clock;
  assign axi_reset = reset;
  assign axi_io_arready = axi_mem_arready; // @[TopMain.scala 103:18]
  assign axi_io_rdata = axi_mem_rdata; // @[TopMain.scala 104:16]
  assign axi_io_icache_rdata = axi_mem_icache_rdata; // @[TopMain.scala 105:23]
  assign axi_io_rvalid = axi_mem_rvalid; // @[TopMain.scala 106:17]
  assign axi_io_awready = axi_mem_awready; // @[TopMain.scala 108:18]
  assign axi_io_wready = axi_mem_wready; // @[TopMain.scala 109:17]
  assign axi_io_bvalid = axi_mem_bvalid; // @[TopMain.scala 110:17]
  assign axi_io_inst_sram_req = icache_io_rd_req; // @[TopMain.scala 95:24]
  assign axi_io_inst_sram_addr = {{32'd0}, icache_io_rd_addr}; // @[TopMain.scala 97:25]
  assign axi_io_data_sram_req = mem_io_data_sram_req; // @[TopMain.scala 98:24]
  assign axi_io_data_sram_wr = mem_io_data_sram_we; // @[TopMain.scala 99:23]
  assign axi_io_data_sram_wstrb = mem_io_data_sram_wmask; // @[TopMain.scala 102:26]
  assign axi_io_data_sram_addr = {{32'd0}, mem_io_data_sram_addr}; // @[TopMain.scala 100:25]
  assign axi_io_data_sram_wdata = mem_io_data_sram_wdata; // @[TopMain.scala 101:26]
  assign axi_mem_reset = reset; // @[TopMain.scala 127:20]
  assign axi_mem_clock = clock; // @[TopMain.scala 128:20]
  assign axi_mem_arid = axi_io_arid; // @[TopMain.scala 129:19]
  assign axi_mem_araddr = axi_io_araddr; // @[TopMain.scala 130:21]
  assign axi_mem_arvalid = axi_io_arvalid; // @[TopMain.scala 131:22]
  assign axi_mem_rready = axi_io_rready; // @[TopMain.scala 133:21]
  assign axi_mem_awid = 4'h1; // @[TopMain.scala 135:19]
  assign axi_mem_awaddr = axi_io_awaddr; // @[TopMain.scala 136:21]
  assign axi_mem_awvalid = axi_io_awvalid; // @[TopMain.scala 137:22]
  assign axi_mem_wdata = axi_io_wdata; // @[TopMain.scala 139:20]
  assign axi_mem_wstrb = axi_io_wstrb; // @[TopMain.scala 140:20]
  assign axi_mem_wvalid = axi_io_wvalid; // @[TopMain.scala 141:21]
  assign axi_mem_bready = axi_io_bready; // @[TopMain.scala 143:21]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_valid = ifu_io_inst_sram_req; // @[TopMain.scala 146:16]
  assign icache_io_addr = ifu_io_inst_sram_addr; // @[TopMain.scala 148:15]
  assign icache_io_rd_rdy = axi_io_inst_sram_addr_ok; // @[TopMain.scala 150:17]
  assign icache_io_rd_data = axi_io_inst_sram_rdata; // @[TopMain.scala 151:18]
  assign icache_io_inst_sram_data_ok = axi_io_inst_sram_data_ok; // @[TopMain.scala 153:28]
endmodule
